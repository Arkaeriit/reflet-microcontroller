module rom01(input clk, input enable, input [6-1:0] addr, output [8-1:0] data);
    reg [8-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            6'h0 : data_reg <= 8'h41;
            6'h1 : data_reg <= 8'h53;
            6'h2 : data_reg <= 8'h52;
            6'h3 : data_reg <= 8'h4D;
            6'h4 : data_reg <= 8'h26;
            6'h5 : data_reg <= 8'h1D;
            6'h6 : data_reg <= 8'h2A;
            6'h7 : data_reg <= 8'h1E;
            6'h8 : data_reg <= 8'h7F;
            6'h9 : data_reg <= 8'h1A;
            6'hA : data_reg <= 8'h28;
            6'hB : data_reg <= 8'h11;
            6'hC : data_reg <= 8'hD1;
            6'hD : data_reg <= 8'h11;
            6'hE : data_reg <= 8'h21;
            6'hF : data_reg <= 8'h31;
            6'h10 : data_reg <= 8'h12;
            6'h11 : data_reg <= 8'h21;
            6'h12 : data_reg <= 8'h32;
            6'h13 : data_reg <= 8'h13;
            6'h14 : data_reg <= 8'h21;
            6'h15 : data_reg <= 8'h33;
            6'h16 : data_reg <= 8'h14;
            6'h17 : data_reg <= 8'h21;
            6'h18 : data_reg <= 8'h34;
            6'h19 : data_reg <= 8'h15;
            6'h1A : data_reg <= 8'h00;
            6'h1B : data_reg <= 8'hD4;
            6'h1C : data_reg <= 8'hC2;
            6'h1D : data_reg <= 8'hD5;
            6'h1E : data_reg <= 8'h41;
            6'h1F : data_reg <= 8'h17;
            6'h20 : data_reg <= 8'hD3;
            6'h21 : data_reg <= 8'h42;
            6'h22 : data_reg <= 8'h18;
            6'h23 : data_reg <= 8'h78;
            6'h24 : data_reg <= 8'h42;
            6'h25 : data_reg <= 8'h57;
            6'h26 : data_reg <= 8'hC3;
            6'h27 : data_reg <= 8'h29;
            6'h28 : data_reg <= 8'h19;
            6'h29 : data_reg <= 8'hD9;
            6'h2A : data_reg <= 8'h1E;
            6'h2B : data_reg <= 8'h00;
            6'h2C : data_reg <= 8'h00;
            6'h2D : data_reg <= 8'hE8;
            default : data_reg <= 0;
        endcase
    assign data = ( enable ? data_reg : 0 );
endmodule
