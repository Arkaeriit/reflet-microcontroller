`define test_instruction_bin_size 828
`define test_instruction_bin 6624'h000e0c2c3d2b3cf04e084c1300993e4e4c123c123d102c3b2d3c0c2c3d2b3cf04e084c1300f33e4e4c123c123d102c3b2d3c0c2c3d2b3cf04e084c1300403e4e4c12003c123d102c3b2d3c3ff02c3d2b3cf04e084c1300383e4e4c123c123d102c3b2d3c0d0c2a311a0e0d0c2a3103f110e1032c3d2b3cf04e084c13ffff3e4e4c123c123d102c3b2d3c314f1809012c3d2b3cf04e084c1302d23e4e4c123c123d102c3b2d3cc11131110c2c3d2b3cf04e084c1302d33e4e4c12003c123d102c3b2d3c0c2a31087c1d3cac103c140c2a310a100b7c103cac153c140c2a31ff10ef7c1a3cac153c143e2c3d2b3cf04e084c1302d23e4e4c123c123d102c3b2d3c092c3d2b3cf04e084c1302543e4e4c123c123d102c3b2d3cd110092c3d2b3cf04e084c1302d23e4e4c123c123d102c3b2d3cd111092c3d2b3cf04e084c1302d23e4e4c123c123d102c3b2d3cc1103e2c3d2b3cf04e084c1302d23e4e4c123c123d102c3b2d3c092c3d2b3cf04e084c1301ee3e4e4c12003c123d102c3b2d3cc11131110c2a31b2160c2a31a21732110c2a31920c2a31831e331d0c2a31727c153cac153c14327c1a3cac1a3c140c2a3162120c2a31627c153cac153c14327c1a3cac1a3c140c2a31527c123cac133c140c2a31527c183cac1c3c14327c143cac163c140c2a31417c1f3cac103c14317c1a3cac103c140c2a3122322c3d2b3cf04e084c130c803e4e4c123c123d102c3b2d3c0c2a31163a2c3d2b3cf04e084c13003a3e4e4c12003c123d102c3b2d3c39f02c3d2b3cf04e084c1300343e4e4c12003c123d102c3b2d3c0d092c3d2b3cf04e084c1300cf3e4e4c123c123d102c3b2d3c01c3223343113141120ff1331032f02c3d2b3cf04e084c1300363e4e4c12003c123d102c3b2d3c31f02c3d2b3cf04e084c1300343e4e4c12003c123d102c3b2d3c0d092c3d2b3cf04e084c1300753e4e4c123c123d102c3b2d3c01c322334311314112e110331032f02c3d2b3cf04e084c1300363e4e4c12003c123d102c3b2d3c31f02c3d2b3cf04e084c1300343e4e4c123c123d102c3b2d3c0d394912e9219000001480003e2c3d2b3cf04e084c1302d83e4e4c123c123d102c3b2d3c3f2c3d2b3cf04e084c13033c3e4e4c123c123d102c3b2d3c4d525341
