//This module is made from the file software/bootloader16.asm
//It is assembled with the macro-assembler and the flags
//-no-prefix, -no-stack-init, -ignore-start and -start-addr 32256
//It is made into a rom with https://github.com/Arkaeriit/ROM_maker

module reflet_bootloader16_rom(input clk, input enable, input [14-1:0] addr, output [15:0] data_out);
    reg [16-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            14'h3F00 : data_reg <= 16'h1003;  //Note: from the CPU's perspective, this is addr 0X7E00
            14'h3F01 : data_reg <= 16'h1432;
            14'h3F02 : data_reg <= 16'h1431;
            14'h3F03 : data_reg <= 16'h103C;
            14'h3F04 : data_reg <= 16'h1F3B;
            14'h3F05 : data_reg <= 16'hAC7B;
            14'h3F06 : data_reg <= 16'h1F3B;
            14'h3F07 : data_reg <= 16'hAC7B;
            14'h3F08 : data_reg <= 16'h103B;
            14'h3F09 : data_reg <= 16'hAC7B;
            14'h3F0A : data_reg <= 16'h103B;
            14'h3F0B : data_reg <= 16'h337B;
            14'h3F0C : data_reg <= 16'h34F3;
            14'h3F0D : data_reg <= 16'h4311;
            14'h3F0E : data_reg <= 16'hF333;
            14'h3F0F : data_reg <= 16'h1F35;
            14'h3F10 : data_reg <= 16'h3343;
            14'h3F11 : data_reg <= 16'h3C14;
            14'h3F12 : data_reg <= 16'h3B10;
            14'h3F13 : data_reg <= 16'h7B10;
            14'h3F14 : data_reg <= 16'h3BAC;
            14'h3F15 : data_reg <= 16'h7B10;
            14'h3F16 : data_reg <= 16'h3BAC;
            14'h3F17 : data_reg <= 16'h7B16;
            14'h3F18 : data_reg <= 16'h3BAC;
            14'h3F19 : data_reg <= 16'h7B13;
            14'h3F1A : data_reg <= 16'h36E3;
            14'h3F1B : data_reg <= 16'h4311;
            14'h3F1C : data_reg <= 16'h2633;
            14'h3F1D : data_reg <= 16'h11E3;
            14'h3F1E : data_reg <= 16'h3343;
            14'h3F1F : data_reg <= 16'hE311;
            14'h3F20 : data_reg <= 16'hC510;
            14'h3F21 : data_reg <= 16'h1401;
            14'h3F22 : data_reg <= 16'h103C;
            14'h3F23 : data_reg <= 16'h173B;
            14'h3F24 : data_reg <= 16'hAC7B;
            14'h3F25 : data_reg <= 16'h1E3B;
            14'h3F26 : data_reg <= 16'hAC7B;
            14'h3F27 : data_reg <= 16'h173B;
            14'h3F28 : data_reg <= 16'hAC7B;
            14'h3F29 : data_reg <= 16'h133B;
            14'h3F2A : data_reg <= 16'h097B;
            14'h3F2B : data_reg <= 16'h4311;
            14'h3F2C : data_reg <= 16'h1133;
            14'h3F2D : data_reg <= 16'h12E3;
            14'h3F2E : data_reg <= 16'h3343;
            14'h3F2F : data_reg <= 16'hE324;
            14'h3F30 : data_reg <= 16'h3C14;
            14'h3F31 : data_reg <= 16'h3B10;
            14'h3F32 : data_reg <= 16'h7B17;
            14'h3F33 : data_reg <= 16'h3BAC;
            14'h3F34 : data_reg <= 16'h7B1E;
            14'h3F35 : data_reg <= 16'h3BAC;
            14'h3F36 : data_reg <= 16'h7B19;
            14'h3F37 : data_reg <= 16'h3BAC;
            14'h3F38 : data_reg <= 16'h7B13;
            14'h3F39 : data_reg <= 16'h113E;
            14'h3F3A : data_reg <= 16'h3343;
            14'h3F3B : data_reg <= 16'hE311;
            14'h3F3C : data_reg <= 16'h4311;
            14'h3F3D : data_reg <= 16'h1433;
            14'h3F3E : data_reg <= 16'h103C;
            14'h3F3F : data_reg <= 16'h103B;
            14'h3F40 : data_reg <= 16'hAC7B;
            14'h3F41 : data_reg <= 16'h103B;
            14'h3F42 : data_reg <= 16'hAC7B;
            14'h3F43 : data_reg <= 16'h1F3B;
            14'h3F44 : data_reg <= 16'hAC7B;
            14'h3F45 : data_reg <= 16'h1F3B;
            14'h3F46 : data_reg <= 16'hE37B;
            14'h3F47 : data_reg <= 16'h4311;
            14'h3F48 : data_reg <= 16'h2533;
            14'h3F49 : data_reg <= 16'h14E3;
            14'h3F4A : data_reg <= 16'h103C;
            14'h3F4B : data_reg <= 16'h1F3B;
            14'h3F4C : data_reg <= 16'hAC7B;
            14'h3F4D : data_reg <= 16'h1F3B;
            14'h3F4E : data_reg <= 16'hAC7B;
            14'h3F4F : data_reg <= 16'h103B;
            14'h3F50 : data_reg <= 16'hAC7B;
            14'h3F51 : data_reg <= 16'h143B;
            14'h3F52 : data_reg <= 16'h337B;
            14'h3F53 : data_reg <= 16'hE31A;
            14'h3F54 : data_reg <= 16'h4311;
            14'h3F55 : data_reg <= 16'h1433;
            14'h3F56 : data_reg <= 16'h103C;
            14'h3F57 : data_reg <= 16'h103B;
            14'h3F58 : data_reg <= 16'hAC7B;
            14'h3F59 : data_reg <= 16'h103B;
            14'h3F5A : data_reg <= 16'hAC7B;
            14'h3F5B : data_reg <= 16'h143B;
            14'h3F5C : data_reg <= 16'hAC7B;
            14'h3F5D : data_reg <= 16'h103B;
            14'h3F5E : data_reg <= 16'hE37B;
            14'h3F5F : data_reg <= 16'h4312;
            14'h3F60 : data_reg <= 16'h1433;
            14'h3F61 : data_reg <= 16'h103C;
            14'h3F62 : data_reg <= 16'h103B;
            14'h3F63 : data_reg <= 16'hAC7B;
            14'h3F64 : data_reg <= 16'h113B;
            14'h3F65 : data_reg <= 16'hAC7B;
            14'h3F66 : data_reg <= 16'h193B;
            14'h3F67 : data_reg <= 16'hAC7B;
            14'h3F68 : data_reg <= 16'h103B;
            14'h3F69 : data_reg <= 16'h367B;
            14'h3F6A : data_reg <= 16'h1431;
            14'h3F6B : data_reg <= 16'h103C;
            14'h3F6C : data_reg <= 16'h1F3B;
            14'h3F6D : data_reg <= 16'hAC7B;
            14'h3F6E : data_reg <= 16'h1F3B;
            14'h3F6F : data_reg <= 16'hAC7B;
            14'h3F70 : data_reg <= 16'h113B;
            14'h3F71 : data_reg <= 16'hAC7B;
            14'h3F72 : data_reg <= 16'h193B;
            14'h3F73 : data_reg <= 16'h377B;
            14'h3F74 : data_reg <= 16'h3C14;
            14'h3F75 : data_reg <= 16'h3B10;
            14'h3F76 : data_reg <= 16'h7B17;
            14'h3F77 : data_reg <= 16'h3BAC;
            14'h3F78 : data_reg <= 16'h7B1F;
            14'h3F79 : data_reg <= 16'h3BAC;
            14'h3F7A : data_reg <= 16'h7B14;
            14'h3F7B : data_reg <= 16'h3BAC;
            14'h3F7C : data_reg <= 16'h7B1E;
            14'h3F7D : data_reg <= 16'h1438;
            14'h3F7E : data_reg <= 16'h103C;
            14'h3F7F : data_reg <= 16'h173B;
            14'h3F80 : data_reg <= 16'hAC7B;
            14'h3F81 : data_reg <= 16'h1F3B;
            14'h3F82 : data_reg <= 16'hAC7B;
            14'h3F83 : data_reg <= 16'h193B;
            14'h3F84 : data_reg <= 16'hAC7B;
            14'h3F85 : data_reg <= 16'h1D3B;
            14'h3F86 : data_reg <= 16'h047B;
            14'h3F87 : data_reg <= 16'h3C14;
            14'h3F88 : data_reg <= 16'h3B10;
            14'h3F89 : data_reg <= 16'h7B17;
            14'h3F8A : data_reg <= 16'h3BAC;
            14'h3F8B : data_reg <= 16'h7B1F;
            14'h3F8C : data_reg <= 16'h3BAC;
            14'h3F8D : data_reg <= 16'h7B1A;
            14'h3F8E : data_reg <= 16'h3BAC;
            14'h3F8F : data_reg <= 16'h7B19;
            14'h3F90 : data_reg <= 16'h1405;
            14'h3F91 : data_reg <= 16'h103C;
            14'h3F92 : data_reg <= 16'h103B;
            14'h3F93 : data_reg <= 16'hAC7B;
            14'h3F94 : data_reg <= 16'h103B;
            14'h3F95 : data_reg <= 16'hAC7B;
            14'h3F96 : data_reg <= 16'h113B;
            14'h3F97 : data_reg <= 16'hAC7B;
            14'h3F98 : data_reg <= 16'h183B;
            14'h3F99 : data_reg <= 16'h3D7B;
            14'h3F9A : data_reg <= 16'h3C14;
            14'h3F9B : data_reg <= 16'h3B10;
            14'h3F9C : data_reg <= 16'h7B17;
            14'h3F9D : data_reg <= 16'h3BAC;
            14'h3F9E : data_reg <= 16'h7B1F;
            14'h3F9F : data_reg <= 16'h3BAC;
            14'h3FA0 : data_reg <= 16'h7B14;
            14'h3FA1 : data_reg <= 16'h3BAC;
            14'h3FA2 : data_reg <= 16'h7B17;
            14'h3FA3 : data_reg <= 16'h003A;
            14'h3FA4 : data_reg <= 16'hC110;
            14'h3FA5 : data_reg <= 16'h0928;
            14'h3FA6 : data_reg <= 16'h3E2A;
            14'h3FA7 : data_reg <= 16'h3D11;
            14'h3FA8 : data_reg <= 16'h3C14;
            14'h3FA9 : data_reg <= 16'h3B10;
            14'h3FAA : data_reg <= 16'h7B1F;
            14'h3FAB : data_reg <= 16'h3BAC;
            14'h3FAC : data_reg <= 16'h7B1F;
            14'h3FAD : data_reg <= 16'h3BAC;
            14'h3FAE : data_reg <= 16'h7B10;
            14'h3FAF : data_reg <= 16'h3BAC;
            14'h3FB0 : data_reg <= 16'h7B14;
            14'h3FB1 : data_reg <= 16'h1031;
            14'h3FB2 : data_reg <= 16'h11E1;
            14'h3FB3 : data_reg <= 16'h3141;
            14'h3FB4 : data_reg <= 16'hE110;
            14'h3FB5 : data_reg <= 16'h4111;
            14'h3FB6 : data_reg <= 16'h1031;
            14'h3FB7 : data_reg <= 16'h19E1;
            14'h3FB8 : data_reg <= 16'h3141;
            14'h3FB9 : data_reg <= 16'hE110;
            14'h3FBA : data_reg <= 16'h4111;
            14'h3FBB : data_reg <= 16'h1031;
            14'h3FBC : data_reg <= 16'h11E1;
            14'h3FBD : data_reg <= 16'h3141;
            14'h3FBE : data_reg <= 16'hE110;
            14'h3FBF : data_reg <= 16'h4111;
            14'h3FC0 : data_reg <= 16'h1031;
            14'h3FC1 : data_reg <= 16'h11E1;
            14'h3FC2 : data_reg <= 16'h3141;
            14'h3FC3 : data_reg <= 16'hE110;
            14'h3FC4 : data_reg <= 16'h4111;
            14'h3FC5 : data_reg <= 16'h1031;
            14'h3FC6 : data_reg <= 16'h31E1;
            14'h3FC7 : data_reg <= 16'h3332;
            14'h3FC8 : data_reg <= 16'h3534;
            14'h3FC9 : data_reg <= 16'h3736;
            14'h3FCA : data_reg <= 16'h3938;
            14'h3FCB : data_reg <= 16'h3B3A;
            14'h3FCC : data_reg <= 16'h3F3C;
            14'h3FCD : data_reg <= 16'h1403;
            14'h3FCE : data_reg <= 16'h343E;
            14'h3FCF : data_reg <= 16'h3126;
            14'h3FD0 : data_reg <= 16'hE310;
            14'h3FD1 : data_reg <= 16'hE2F7;
            14'h3FD2 : data_reg <= 16'h4211;
            14'h3FD3 : data_reg <= 16'h2432;
            14'h3FD4 : data_reg <= 16'h3502;
            14'h3FD5 : data_reg <= 16'hE310;
            14'h3FD6 : data_reg <= 16'h3911;
            14'h3FD7 : data_reg <= 16'h5921;
            14'h3FD8 : data_reg <= 16'h2531;
            14'h3FD9 : data_reg <= 16'h0002;
            default : data_reg <= 0;
        endcase
    assign data_out = ( enable ? data_reg : 0 );
endmodule
