//The cade used to make this rom om is in software/basicInt.asm
module rom3(input clk, input enable, input [7-1:0] addr, output [8-1:0] dataOut);
    reg [8-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            7'h0 : data_reg <= 8'h41;
            7'h1 : data_reg <= 8'h53;
            7'h2 : data_reg <= 8'h52;
            7'h3 : data_reg <= 8'h4D;
            7'h4 : data_reg <= 8'h14;
            7'h5 : data_reg <= 8'h3C;
            7'h6 : data_reg <= 8'h18;
            7'h7 : data_reg <= 8'hAC;
            7'h8 : data_reg <= 8'h3C;
            7'h9 : data_reg <= 8'h14;
            7'hA : data_reg <= 8'h7C;
            7'hB : data_reg <= 8'h31;
            7'hC : data_reg <= 8'h10;
            7'hD : data_reg <= 8'h90;
            7'hE : data_reg <= 8'h32;
            7'hF : data_reg <= 8'hE1;
            7'h10 : data_reg <= 8'h11;
            7'h11 : data_reg <= 8'h41;
            7'h12 : data_reg <= 8'h31;
            7'h13 : data_reg <= 8'h22;
            7'h14 : data_reg <= 8'hE1;
            7'h15 : data_reg <= 8'h11;
            7'h16 : data_reg <= 8'h41;
            7'h17 : data_reg <= 8'h31;
            7'h18 : data_reg <= 8'h22;
            7'h19 : data_reg <= 8'hE1;
            7'h1A : data_reg <= 8'h11;
            7'h1B : data_reg <= 8'h41;
            7'h1C : data_reg <= 8'h31;
            7'h1D : data_reg <= 8'h22;
            7'h1E : data_reg <= 8'hE1;
            7'h1F : data_reg <= 8'h11;
            7'h20 : data_reg <= 8'h41;
            7'h21 : data_reg <= 8'h31;
            7'h22 : data_reg <= 8'h11;
            7'h23 : data_reg <= 8'hE1;
            7'h24 : data_reg <= 8'h41;
            7'h25 : data_reg <= 8'h31;
            7'h26 : data_reg <= 8'h12;
            7'h27 : data_reg <= 8'hE1;
            7'h28 : data_reg <= 8'h11;
            7'h29 : data_reg <= 8'h41;
            7'h2A : data_reg <= 8'h31;
            7'h2B : data_reg <= 8'h11;
            7'h2C : data_reg <= 8'h41;
            7'h2D : data_reg <= 8'h31;
            7'h2E : data_reg <= 8'h3C;
            7'h2F : data_reg <= 8'h2D;
            7'h30 : data_reg <= 8'h3B;
            7'h31 : data_reg <= 8'h2C;
            7'h32 : data_reg <= 8'h10;
            7'h33 : data_reg <= 8'h3D;
            7'h34 : data_reg <= 8'h11;
            7'h35 : data_reg <= 8'h3C;
            7'h36 : data_reg <= 8'h00;
            7'h37 : data_reg <= 8'h00;
            7'h38 : data_reg <= 8'h00;
            7'h39 : data_reg <= 8'h00;
            7'h3A : data_reg <= 8'h12;
            7'h3B : data_reg <= 8'h4C;
            7'h3C : data_reg <= 8'h4E;
            7'h3D : data_reg <= 8'h3E;
            7'h3E : data_reg <= 8'h6F;
            7'h3F : data_reg <= 8'h13;
            7'h40 : data_reg <= 8'h4C;
            7'h41 : data_reg <= 8'h08;
            7'h42 : data_reg <= 8'h4E;
            7'h43 : data_reg <= 8'hF0;
            7'h44 : data_reg <= 8'h3C;
            7'h45 : data_reg <= 8'h2B;
            7'h46 : data_reg <= 8'h3D;
            7'h47 : data_reg <= 8'h2C;
            7'h48 : data_reg <= 8'h06;
            7'h49 : data_reg <= 8'h14;
            7'h4A : data_reg <= 8'h3C;
            7'h4B : data_reg <= 8'h12;
            7'h4C : data_reg <= 8'hAC;
            7'h4D : data_reg <= 8'h3C;
            7'h4E : data_reg <= 8'h10;
            7'h4F : data_reg <= 8'h7C;
            7'h50 : data_reg <= 8'h3D;
            7'h51 : data_reg <= 8'h3C;
            7'h52 : data_reg <= 8'h2D;
            7'h53 : data_reg <= 8'h3B;
            7'h54 : data_reg <= 8'h2C;
            7'h55 : data_reg <= 8'h10;
            7'h56 : data_reg <= 8'h3D;
            7'h57 : data_reg <= 8'h11;
            7'h58 : data_reg <= 8'h3C;
            7'h59 : data_reg <= 8'h00;
            7'h5A : data_reg <= 8'h00;
            7'h5B : data_reg <= 8'h00;
            7'h5C : data_reg <= 8'h00;
            7'h5D : data_reg <= 8'h12;
            7'h5E : data_reg <= 8'h4C;
            7'h5F : data_reg <= 8'h4E;
            7'h60 : data_reg <= 8'h3E;
            7'h61 : data_reg <= 8'h6B;
            7'h62 : data_reg <= 8'h13;
            7'h63 : data_reg <= 8'h4C;
            7'h64 : data_reg <= 8'h08;
            7'h65 : data_reg <= 8'h4E;
            7'h66 : data_reg <= 8'hF0;
            7'h67 : data_reg <= 8'h3C;
            7'h68 : data_reg <= 8'h2B;
            7'h69 : data_reg <= 8'h3D;
            7'h6A : data_reg <= 8'h2C;
            7'h6B : data_reg <= 8'h00;
            7'h6C : data_reg <= 8'h00;
            7'h6D : data_reg <= 8'h3E;
            7'h6E : data_reg <= 8'h0E;
            7'h6F : data_reg <= 8'h32;
            7'h70 : data_reg <= 8'h0F;
            7'h71 : data_reg <= 8'h10;
            7'h72 : data_reg <= 8'hE1;
            7'h73 : data_reg <= 8'h22;
            7'h74 : data_reg <= 8'h02;
            default : data_reg <= 0;
        endcase
    assign dataOut = ( enable ? data_reg : 0 );
endmodule
