module rom07(input clk, input enable, input [14-1:0] addr, output [16-1:0] data);
    reg [16-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            14'h0 : data_reg <= 16'h5341;
            14'h1 : data_reg <= 16'h4D52;
            14'h2 : data_reg <= 16'h1C28;
            14'h3 : data_reg <= 16'h8C22;
            14'h4 : data_reg <= 16'h9C6D;
            14'h5 : data_reg <= 16'h6D8C;
            14'h6 : data_reg <= 16'h0D1D;
            14'h7 : data_reg <= 16'h281B;
            14'h8 : data_reg <= 16'h221C;
            14'h9 : data_reg <= 16'h6D8C;
            14'hA : data_reg <= 16'h8C9C;
            14'hB : data_reg <= 16'h1D6D;
            14'hC : data_reg <= 16'h1C22;
            14'hD : data_reg <= 16'h3C22;
            14'hE : data_reg <= 16'h1E3E;
            14'hF : data_reg <= 16'h8000;
            14'h10 : data_reg <= 16'h3C23;
            14'h11 : data_reg <= 16'h3EE5;
            14'h12 : data_reg <= 16'h1CD0;
            14'h13 : data_reg <= 16'h1D0B;
            14'h14 : data_reg <= 16'h1F0C;
            14'h15 : data_reg <= 16'h1B0D;
            14'h16 : data_reg <= 16'h1C28;
            14'h17 : data_reg <= 16'h8C22;
            14'h18 : data_reg <= 16'h9C6D;
            14'h19 : data_reg <= 16'h6D8C;
            14'h1A : data_reg <= 16'h221D;
            14'h1B : data_reg <= 16'h001C;
            14'h1C : data_reg <= 16'h3C22;
            14'h1D : data_reg <= 16'h1E3E;
            14'h1E : data_reg <= 16'h01C9;
            14'h1F : data_reg <= 16'h3C23;
            14'h20 : data_reg <= 16'h3EE5;
            14'h21 : data_reg <= 16'h1CD0;
            14'h22 : data_reg <= 16'h1D0B;
            14'h23 : data_reg <= 16'h1E0C;
            14'h24 : data_reg <= 16'h7D00;
            14'h25 : data_reg <= 16'h8000;
            14'h26 : data_reg <= 16'hFF00;
            14'h27 : data_reg <= 16'hFF04;
            14'h28 : data_reg <= 16'hFF08;
            14'h29 : data_reg <= 16'hFF10;
            14'h2A : data_reg <= 16'hFF13;
            14'h2B : data_reg <= 16'hFF16;
            14'h2C : data_reg <= 16'hFF1A;
            14'h2D : data_reg <= 16'hFF1C;
            14'h2E : data_reg <= 16'hFF1F;
            14'h2F : data_reg <= 16'hFF21;
            14'h30 : data_reg <= 16'hFF22;
            14'h31 : data_reg <= 16'h021C;
            14'h32 : data_reg <= 16'h0CE4;
            14'h33 : data_reg <= 16'h041C;
            14'h34 : data_reg <= 16'h0CE4;
            14'h35 : data_reg <= 16'h1B0D;
            14'h36 : data_reg <= 16'h1C28;
            14'h37 : data_reg <= 16'h8C22;
            14'h38 : data_reg <= 16'h9C6D;
            14'h39 : data_reg <= 16'h6D8C;
            14'h3A : data_reg <= 16'h221D;
            14'h3B : data_reg <= 16'h001C;
            14'h3C : data_reg <= 16'h3C22;
            14'h3D : data_reg <= 16'h1E3E;
            14'h3E : data_reg <= 16'h0056;
            14'h3F : data_reg <= 16'h3C23;
            14'h40 : data_reg <= 16'h3EE5;
            14'h41 : data_reg <= 16'h1CD0;
            14'h42 : data_reg <= 16'h1D0B;
            14'h43 : data_reg <= 16'hD00C;
            14'h44 : data_reg <= 16'h0D12;
            14'h45 : data_reg <= 16'h281B;
            14'h46 : data_reg <= 16'h221C;
            14'h47 : data_reg <= 16'h6D8C;
            14'h48 : data_reg <= 16'h8C9C;
            14'h49 : data_reg <= 16'h1D6D;
            14'h4A : data_reg <= 16'h1C22;
            14'h4B : data_reg <= 16'h3C22;
            14'h4C : data_reg <= 16'h1E3E;
            14'h4D : data_reg <= 16'h00A6;
            14'h4E : data_reg <= 16'h3C23;
            14'h4F : data_reg <= 16'h3EE5;
            14'h50 : data_reg <= 16'h1CD0;
            14'h51 : data_reg <= 16'h1D0B;
            14'h52 : data_reg <= 16'h140C;
            14'h53 : data_reg <= 16'h1B0D;
            14'h54 : data_reg <= 16'h1C28;
            14'h55 : data_reg <= 16'h8C21;
            14'h56 : data_reg <= 16'h9C6D;
            14'h57 : data_reg <= 16'h6D8C;
            14'h58 : data_reg <= 16'hD21D;
            14'h59 : data_reg <= 16'h0B1C;
            14'h5A : data_reg <= 16'h0C1D;
            14'h5B : data_reg <= 16'h201C;
            14'h5C : data_reg <= 16'h04AC;
            14'h5D : data_reg <= 16'h21E0;
            14'h5E : data_reg <= 16'h1432;
            14'h5F : data_reg <= 16'h1B01;
            14'h60 : data_reg <= 16'h1C28;
            14'h61 : data_reg <= 16'h8C21;
            14'h62 : data_reg <= 16'h9C6D;
            14'h63 : data_reg <= 16'h6D8C;
            14'h64 : data_reg <= 16'h1C6D;
            14'h65 : data_reg <= 16'h6C0D;
            14'h66 : data_reg <= 16'h0B1D;
            14'h67 : data_reg <= 16'h1BC4;
            14'h68 : data_reg <= 16'h6D0C;
            14'h69 : data_reg <= 16'h0B1D;
            14'h6A : data_reg <= 16'h1B20;
            14'h6B : data_reg <= 16'h1C28;
            14'h6C : data_reg <= 16'h8C21;
            14'h6D : data_reg <= 16'h9C6D;
            14'h6E : data_reg <= 16'h6D8C;
            14'h6F : data_reg <= 16'h1C6D;
            14'h70 : data_reg <= 16'h6C0D;
            14'h71 : data_reg <= 16'h0B1D;
            14'h72 : data_reg <= 16'h1BC2;
            14'h73 : data_reg <= 16'h6D0C;
            14'h74 : data_reg <= 16'h0B1D;
            14'h75 : data_reg <= 16'hE31C;
            14'h76 : data_reg <= 16'h0C14;
            14'h77 : data_reg <= 16'hE31C;
            14'h78 : data_reg <= 16'h0C12;
            14'h79 : data_reg <= 16'h1CE2;
            14'h7A : data_reg <= 16'hE401;
            14'h7B : data_reg <= 16'h2A0C;
            14'h7C : data_reg <= 16'h0D11;
            14'h7D : data_reg <= 16'h281B;
            14'h7E : data_reg <= 16'h221C;
            14'h7F : data_reg <= 16'h6D8C;
            14'h80 : data_reg <= 16'h8C9C;
            14'h81 : data_reg <= 16'h1D6D;
            14'h82 : data_reg <= 16'h1C22;
            14'h83 : data_reg <= 16'h3C22;
            14'h84 : data_reg <= 16'h1E3E;
            14'h85 : data_reg <= 16'h0062;
            14'h86 : data_reg <= 16'h3C23;
            14'h87 : data_reg <= 16'h3EE5;
            14'h88 : data_reg <= 16'h1CD0;
            14'h89 : data_reg <= 16'h1D0B;
            14'h8A : data_reg <= 16'hE10C;
            14'h8B : data_reg <= 16'h112D;
            14'h8C : data_reg <= 16'h1B0D;
            14'h8D : data_reg <= 16'h1C28;
            14'h8E : data_reg <= 16'h8C22;
            14'h8F : data_reg <= 16'h9C6D;
            14'h90 : data_reg <= 16'h6D8C;
            14'h91 : data_reg <= 16'h221D;
            14'h92 : data_reg <= 16'h001C;
            14'h93 : data_reg <= 16'h3C22;
            14'h94 : data_reg <= 16'h1E3E;
            14'h95 : data_reg <= 16'h0062;
            14'h96 : data_reg <= 16'h3C23;
            14'h97 : data_reg <= 16'h3EE5;
            14'h98 : data_reg <= 16'h1CD0;
            14'h99 : data_reg <= 16'h1D0B;
            14'h9A : data_reg <= 16'hE10C;
            14'h9B : data_reg <= 16'hE31C;
            14'h9C : data_reg <= 16'h0C11;
            14'h9D : data_reg <= 16'h1CE2;
            14'h9E : data_reg <= 16'hE402;
            14'h9F : data_reg <= 16'h1C0C;
            14'hA0 : data_reg <= 16'hE403;
            14'hA1 : data_reg <= 16'h0D0C;
            14'hA2 : data_reg <= 16'h281B;
            14'hA3 : data_reg <= 16'h221C;
            14'hA4 : data_reg <= 16'h6D8C;
            14'hA5 : data_reg <= 16'h8C9C;
            14'hA6 : data_reg <= 16'h1D6D;
            14'hA7 : data_reg <= 16'h1C22;
            14'hA8 : data_reg <= 16'h3C22;
            14'hA9 : data_reg <= 16'h1E3E;
            14'hAA : data_reg <= 16'h0056;
            14'hAB : data_reg <= 16'h3C23;
            14'hAC : data_reg <= 16'h3EE5;
            14'hAD : data_reg <= 16'h1CD0;
            14'hAE : data_reg <= 16'h1D0B;
            14'hAF : data_reg <= 16'hD00C;
            14'hB0 : data_reg <= 16'h2212;
            14'hB1 : data_reg <= 16'h1232;
            14'hB2 : data_reg <= 16'h1B0D;
            14'hB3 : data_reg <= 16'h1C28;
            14'hB4 : data_reg <= 16'h8C22;
            14'hB5 : data_reg <= 16'h9C6D;
            14'hB6 : data_reg <= 16'h6D8C;
            14'hB7 : data_reg <= 16'h221D;
            14'hB8 : data_reg <= 16'h001C;
            14'hB9 : data_reg <= 16'h3C22;
            14'hBA : data_reg <= 16'h1E3E;
            14'hBB : data_reg <= 16'h0199;
            14'hBC : data_reg <= 16'h3C23;
            14'hBD : data_reg <= 16'h3EE5;
            14'hBE : data_reg <= 16'h1CD0;
            14'hBF : data_reg <= 16'h1D0B;
            14'hC0 : data_reg <= 16'h130C;
            14'hC1 : data_reg <= 16'h1B21;
            14'hC2 : data_reg <= 16'h1C28;
            14'hC3 : data_reg <= 16'h8C21;
            14'hC4 : data_reg <= 16'h9C6D;
            14'hC5 : data_reg <= 16'h6D8C;
            14'hC6 : data_reg <= 16'h1C6D;
            14'hC7 : data_reg <= 16'h6C0D;
            14'hC8 : data_reg <= 16'h0B1D;
            14'hC9 : data_reg <= 16'h1BC2;
            14'hCA : data_reg <= 16'h6D0C;
            14'hCB : data_reg <= 16'h0B1D;
            14'hCC : data_reg <= 16'h0D11;
            14'hCD : data_reg <= 16'h281B;
            14'hCE : data_reg <= 16'h211C;
            14'hCF : data_reg <= 16'h6D8C;
            14'hD0 : data_reg <= 16'h8C9C;
            14'hD1 : data_reg <= 16'h1D6D;
            14'hD2 : data_reg <= 16'h1CD2;
            14'hD3 : data_reg <= 16'h1D0B;
            14'hD4 : data_reg <= 16'hA10C;
            14'hD5 : data_reg <= 16'hE003;
            14'hD6 : data_reg <= 16'h3221;
            14'hD7 : data_reg <= 16'h0D12;
            14'hD8 : data_reg <= 16'h281B;
            14'hD9 : data_reg <= 16'h211C;
            14'hDA : data_reg <= 16'h6D8C;
            14'hDB : data_reg <= 16'h8C9C;
            14'hDC : data_reg <= 16'h1D6D;
            14'hDD : data_reg <= 16'h1CD2;
            14'hDE : data_reg <= 16'h1D0B;
            14'hDF : data_reg <= 16'h110C;
            14'hE0 : data_reg <= 16'hE31C;
            14'hE1 : data_reg <= 16'h0C13;
            14'hE2 : data_reg <= 16'hE31C;
            14'hE3 : data_reg <= 16'h0C12;
            14'hE4 : data_reg <= 16'h0DE2;
            14'hE5 : data_reg <= 16'h281B;
            14'hE6 : data_reg <= 16'h221C;
            14'hE7 : data_reg <= 16'h6D8C;
            14'hE8 : data_reg <= 16'h8C9C;
            14'hE9 : data_reg <= 16'h1D6D;
            14'hEA : data_reg <= 16'h1C22;
            14'hEB : data_reg <= 16'h3C22;
            14'hEC : data_reg <= 16'h1E3E;
            14'hED : data_reg <= 16'h013B;
            14'hEE : data_reg <= 16'h3C23;
            14'hEF : data_reg <= 16'h3EE5;
            14'hF0 : data_reg <= 16'h1CD0;
            14'hF1 : data_reg <= 16'h1D0B;
            14'hF2 : data_reg <= 16'hE10C;
            14'hF3 : data_reg <= 16'h1B0D;
            14'hF4 : data_reg <= 16'h1C28;
            14'hF5 : data_reg <= 16'h8C22;
            14'hF6 : data_reg <= 16'h9C6D;
            14'hF7 : data_reg <= 16'h6D8C;
            14'hF8 : data_reg <= 16'h221D;
            14'hF9 : data_reg <= 16'h001C;
            14'hFA : data_reg <= 16'h3C22;
            14'hFB : data_reg <= 16'h1E3E;
            14'hFC : data_reg <= 16'h0062;
            14'hFD : data_reg <= 16'h3C23;
            14'hFE : data_reg <= 16'h3EE5;
            14'hFF : data_reg <= 16'h1CD0;
            14'h100 : data_reg <= 16'h1D0B;
            14'h101 : data_reg <= 16'hE10C;
            14'h102 : data_reg <= 16'h1B0D;
            14'h103 : data_reg <= 16'h1C28;
            14'h104 : data_reg <= 16'h8C22;
            14'h105 : data_reg <= 16'h9C6D;
            14'h106 : data_reg <= 16'h6D8C;
            14'h107 : data_reg <= 16'h221D;
            14'h108 : data_reg <= 16'h001C;
            14'h109 : data_reg <= 16'h3C22;
            14'h10A : data_reg <= 16'h1E3E;
            14'h10B : data_reg <= 16'h01C9;
            14'h10C : data_reg <= 16'h3C23;
            14'h10D : data_reg <= 16'h3EE5;
            14'h10E : data_reg <= 16'h1CD0;
            14'h10F : data_reg <= 16'h1D0B;
            14'h110 : data_reg <= 16'h1E0C;
            default : data_reg <= 0;
        endcase
    assign data = ( enable ? data_reg : 0 );
endmodule
