//This module is made from the file software/bootloader16.rasm
//It is assembled with the macro-assembler and the flags
//-no-prefix, -no-stack-init, -ignore-start and -start-addr 32256
module reflet_bootloader16_rom(input clk, input enable, input [14:0] addr, output [7:0] data_out);
reg [7:0] ret; assign data_out = (enable ? ret : 8'h0);
always @ (posedge clk)
case(addr)
  15'h7e00 : ret = 8'h10;
  15'h7e01 : ret = 8'h32;
  15'h7e02 : ret = 8'h14;
  15'h7e03 : ret = 8'h31;
  15'h7e04 : ret = 8'h14;
  15'h7e05 : ret = 8'h3c;
  15'h7e06 : ret = 8'h10;
  15'h7e07 : ret = 8'h3b;
  15'h7e08 : ret = 8'h1f;
  15'h7e09 : ret = 8'h7b;
  15'h7e0a : ret = 8'hac;
  15'h7e0b : ret = 8'h3b;
  15'h7e0c : ret = 8'h1f;
  15'h7e0d : ret = 8'h7b;
  15'h7e0e : ret = 8'hac;
  15'h7e0f : ret = 8'h3b;
  15'h7e10 : ret = 8'h10;
  15'h7e11 : ret = 8'h7b;
  15'h7e12 : ret = 8'hac;
  15'h7e13 : ret = 8'h3b;
  15'h7e14 : ret = 8'h10;
  15'h7e15 : ret = 8'h7b;
  15'h7e16 : ret = 8'h33;
  15'h7e17 : ret = 8'hf3;
  15'h7e18 : ret = 8'h34;
  15'h7e19 : ret = 8'h11;
  15'h7e1a : ret = 8'h43;
  15'h7e1b : ret = 8'h33;
  15'h7e1c : ret = 8'hf3;
  15'h7e1d : ret = 8'h35;
  15'h7e1e : ret = 8'h1f;
  15'h7e1f : ret = 8'h43;
  15'h7e20 : ret = 8'h33;
  15'h7e21 : ret = 8'h14;
  15'h7e22 : ret = 8'h3c;
  15'h7e23 : ret = 8'h10;
  15'h7e24 : ret = 8'h3b;
  15'h7e25 : ret = 8'h10;
  15'h7e26 : ret = 8'h7b;
  15'h7e27 : ret = 8'hac;
  15'h7e28 : ret = 8'h3b;
  15'h7e29 : ret = 8'h10;
  15'h7e2a : ret = 8'h7b;
  15'h7e2b : ret = 8'hac;
  15'h7e2c : ret = 8'h3b;
  15'h7e2d : ret = 8'h16;
  15'h7e2e : ret = 8'h7b;
  15'h7e2f : ret = 8'hac;
  15'h7e30 : ret = 8'h3b;
  15'h7e31 : ret = 8'h13;
  15'h7e32 : ret = 8'h7b;
  15'h7e33 : ret = 8'he3;
  15'h7e34 : ret = 8'h36;
  15'h7e35 : ret = 8'h11;
  15'h7e36 : ret = 8'h43;
  15'h7e37 : ret = 8'h33;
  15'h7e38 : ret = 8'h26;
  15'h7e39 : ret = 8'he3;
  15'h7e3a : ret = 8'h11;
  15'h7e3b : ret = 8'h43;
  15'h7e3c : ret = 8'h33;
  15'h7e3d : ret = 8'h11;
  15'h7e3e : ret = 8'he3;
  15'h7e3f : ret = 8'h10;
  15'h7e40 : ret = 8'hc5;
  15'h7e41 : ret = 8'h1;
  15'h7e42 : ret = 8'h14;
  15'h7e43 : ret = 8'h3c;
  15'h7e44 : ret = 8'h10;
  15'h7e45 : ret = 8'h3b;
  15'h7e46 : ret = 8'h17;
  15'h7e47 : ret = 8'h7b;
  15'h7e48 : ret = 8'hac;
  15'h7e49 : ret = 8'h3b;
  15'h7e4a : ret = 8'h1e;
  15'h7e4b : ret = 8'h7b;
  15'h7e4c : ret = 8'hac;
  15'h7e4d : ret = 8'h3b;
  15'h7e4e : ret = 8'h17;
  15'h7e4f : ret = 8'h7b;
  15'h7e50 : ret = 8'hac;
  15'h7e51 : ret = 8'h3b;
  15'h7e52 : ret = 8'h12;
  15'h7e53 : ret = 8'h7b;
  15'h7e54 : ret = 8'h9;
  15'h7e55 : ret = 8'h11;
  15'h7e56 : ret = 8'h43;
  15'h7e57 : ret = 8'h33;
  15'h7e58 : ret = 8'h11;
  15'h7e59 : ret = 8'he3;
  15'h7e5a : ret = 8'h12;
  15'h7e5b : ret = 8'h43;
  15'h7e5c : ret = 8'h33;
  15'h7e5d : ret = 8'h24;
  15'h7e5e : ret = 8'he3;
  15'h7e5f : ret = 8'h14;
  15'h7e60 : ret = 8'h3c;
  15'h7e61 : ret = 8'h10;
  15'h7e62 : ret = 8'h3b;
  15'h7e63 : ret = 8'h17;
  15'h7e64 : ret = 8'h7b;
  15'h7e65 : ret = 8'hac;
  15'h7e66 : ret = 8'h3b;
  15'h7e67 : ret = 8'h1e;
  15'h7e68 : ret = 8'h7b;
  15'h7e69 : ret = 8'hac;
  15'h7e6a : ret = 8'h3b;
  15'h7e6b : ret = 8'h19;
  15'h7e6c : ret = 8'h7b;
  15'h7e6d : ret = 8'hac;
  15'h7e6e : ret = 8'h3b;
  15'h7e6f : ret = 8'h12;
  15'h7e70 : ret = 8'h7b;
  15'h7e71 : ret = 8'h8;
  15'h7e72 : ret = 8'h11;
  15'h7e73 : ret = 8'h43;
  15'h7e74 : ret = 8'h33;
  15'h7e75 : ret = 8'h11;
  15'h7e76 : ret = 8'he3;
  15'h7e77 : ret = 8'h11;
  15'h7e78 : ret = 8'h43;
  15'h7e79 : ret = 8'h33;
  15'h7e7a : ret = 8'h14;
  15'h7e7b : ret = 8'h3c;
  15'h7e7c : ret = 8'h10;
  15'h7e7d : ret = 8'h3b;
  15'h7e7e : ret = 8'h10;
  15'h7e7f : ret = 8'h7b;
  15'h7e80 : ret = 8'hac;
  15'h7e81 : ret = 8'h3b;
  15'h7e82 : ret = 8'h10;
  15'h7e83 : ret = 8'h7b;
  15'h7e84 : ret = 8'hac;
  15'h7e85 : ret = 8'h3b;
  15'h7e86 : ret = 8'h1f;
  15'h7e87 : ret = 8'h7b;
  15'h7e88 : ret = 8'hac;
  15'h7e89 : ret = 8'h3b;
  15'h7e8a : ret = 8'h1f;
  15'h7e8b : ret = 8'h7b;
  15'h7e8c : ret = 8'he3;
  15'h7e8d : ret = 8'h11;
  15'h7e8e : ret = 8'h43;
  15'h7e8f : ret = 8'h33;
  15'h7e90 : ret = 8'h25;
  15'h7e91 : ret = 8'he3;
  15'h7e92 : ret = 8'h14;
  15'h7e93 : ret = 8'h3c;
  15'h7e94 : ret = 8'h10;
  15'h7e95 : ret = 8'h3b;
  15'h7e96 : ret = 8'h1f;
  15'h7e97 : ret = 8'h7b;
  15'h7e98 : ret = 8'hac;
  15'h7e99 : ret = 8'h3b;
  15'h7e9a : ret = 8'h1f;
  15'h7e9b : ret = 8'h7b;
  15'h7e9c : ret = 8'hac;
  15'h7e9d : ret = 8'h3b;
  15'h7e9e : ret = 8'h10;
  15'h7e9f : ret = 8'h7b;
  15'h7ea0 : ret = 8'hac;
  15'h7ea1 : ret = 8'h3b;
  15'h7ea2 : ret = 8'h14;
  15'h7ea3 : ret = 8'h7b;
  15'h7ea4 : ret = 8'h33;
  15'h7ea5 : ret = 8'h1a;
  15'h7ea6 : ret = 8'he3;
  15'h7ea7 : ret = 8'h11;
  15'h7ea8 : ret = 8'h43;
  15'h7ea9 : ret = 8'h33;
  15'h7eaa : ret = 8'h14;
  15'h7eab : ret = 8'h3c;
  15'h7eac : ret = 8'h10;
  15'h7ead : ret = 8'h3b;
  15'h7eae : ret = 8'h10;
  15'h7eaf : ret = 8'h7b;
  15'h7eb0 : ret = 8'hac;
  15'h7eb1 : ret = 8'h3b;
  15'h7eb2 : ret = 8'h10;
  15'h7eb3 : ret = 8'h7b;
  15'h7eb4 : ret = 8'hac;
  15'h7eb5 : ret = 8'h3b;
  15'h7eb6 : ret = 8'h14;
  15'h7eb7 : ret = 8'h7b;
  15'h7eb8 : ret = 8'hac;
  15'h7eb9 : ret = 8'h3b;
  15'h7eba : ret = 8'h10;
  15'h7ebb : ret = 8'h7b;
  15'h7ebc : ret = 8'he3;
  15'h7ebd : ret = 8'h12;
  15'h7ebe : ret = 8'h43;
  15'h7ebf : ret = 8'h33;
  15'h7ec0 : ret = 8'h14;
  15'h7ec1 : ret = 8'h3c;
  15'h7ec2 : ret = 8'h10;
  15'h7ec3 : ret = 8'h3b;
  15'h7ec4 : ret = 8'h10;
  15'h7ec5 : ret = 8'h7b;
  15'h7ec6 : ret = 8'hac;
  15'h7ec7 : ret = 8'h3b;
  15'h7ec8 : ret = 8'h11;
  15'h7ec9 : ret = 8'h7b;
  15'h7eca : ret = 8'hac;
  15'h7ecb : ret = 8'h3b;
  15'h7ecc : ret = 8'h19;
  15'h7ecd : ret = 8'h7b;
  15'h7ece : ret = 8'hac;
  15'h7ecf : ret = 8'h3b;
  15'h7ed0 : ret = 8'h10;
  15'h7ed1 : ret = 8'h7b;
  15'h7ed2 : ret = 8'h36;
  15'h7ed3 : ret = 8'h31;
  15'h7ed4 : ret = 8'h14;
  15'h7ed5 : ret = 8'h3c;
  15'h7ed6 : ret = 8'h10;
  15'h7ed7 : ret = 8'h3b;
  15'h7ed8 : ret = 8'h1f;
  15'h7ed9 : ret = 8'h7b;
  15'h7eda : ret = 8'hac;
  15'h7edb : ret = 8'h3b;
  15'h7edc : ret = 8'h1f;
  15'h7edd : ret = 8'h7b;
  15'h7ede : ret = 8'hac;
  15'h7edf : ret = 8'h3b;
  15'h7ee0 : ret = 8'h11;
  15'h7ee1 : ret = 8'h7b;
  15'h7ee2 : ret = 8'hac;
  15'h7ee3 : ret = 8'h3b;
  15'h7ee4 : ret = 8'h19;
  15'h7ee5 : ret = 8'h7b;
  15'h7ee6 : ret = 8'h37;
  15'h7ee7 : ret = 8'h14;
  15'h7ee8 : ret = 8'h3c;
  15'h7ee9 : ret = 8'h10;
  15'h7eea : ret = 8'h3b;
  15'h7eeb : ret = 8'h17;
  15'h7eec : ret = 8'h7b;
  15'h7eed : ret = 8'hac;
  15'h7eee : ret = 8'h3b;
  15'h7eef : ret = 8'h1f;
  15'h7ef0 : ret = 8'h7b;
  15'h7ef1 : ret = 8'hac;
  15'h7ef2 : ret = 8'h3b;
  15'h7ef3 : ret = 8'h14;
  15'h7ef4 : ret = 8'h7b;
  15'h7ef5 : ret = 8'hac;
  15'h7ef6 : ret = 8'h3b;
  15'h7ef7 : ret = 8'h1d;
  15'h7ef8 : ret = 8'h7b;
  15'h7ef9 : ret = 8'h38;
  15'h7efa : ret = 8'h14;
  15'h7efb : ret = 8'h3c;
  15'h7efc : ret = 8'h10;
  15'h7efd : ret = 8'h3b;
  15'h7efe : ret = 8'h17;
  15'h7eff : ret = 8'h7b;
  15'h7f00 : ret = 8'hac;
  15'h7f01 : ret = 8'h3b;
  15'h7f02 : ret = 8'h1f;
  15'h7f03 : ret = 8'h7b;
  15'h7f04 : ret = 8'hac;
  15'h7f05 : ret = 8'h3b;
  15'h7f06 : ret = 8'h19;
  15'h7f07 : ret = 8'h7b;
  15'h7f08 : ret = 8'hac;
  15'h7f09 : ret = 8'h3b;
  15'h7f0a : ret = 8'h1b;
  15'h7f0b : ret = 8'h7b;
  15'h7f0c : ret = 8'h4;
  15'h7f0d : ret = 8'h14;
  15'h7f0e : ret = 8'h3c;
  15'h7f0f : ret = 8'h10;
  15'h7f10 : ret = 8'h3b;
  15'h7f11 : ret = 8'h17;
  15'h7f12 : ret = 8'h7b;
  15'h7f13 : ret = 8'hac;
  15'h7f14 : ret = 8'h3b;
  15'h7f15 : ret = 8'h1f;
  15'h7f16 : ret = 8'h7b;
  15'h7f17 : ret = 8'hac;
  15'h7f18 : ret = 8'h3b;
  15'h7f19 : ret = 8'h1a;
  15'h7f1a : ret = 8'h7b;
  15'h7f1b : ret = 8'hac;
  15'h7f1c : ret = 8'h3b;
  15'h7f1d : ret = 8'h17;
  15'h7f1e : ret = 8'h7b;
  15'h7f1f : ret = 8'h5;
  15'h7f20 : ret = 8'h14;
  15'h7f21 : ret = 8'h3c;
  15'h7f22 : ret = 8'h10;
  15'h7f23 : ret = 8'h3b;
  15'h7f24 : ret = 8'h10;
  15'h7f25 : ret = 8'h7b;
  15'h7f26 : ret = 8'hac;
  15'h7f27 : ret = 8'h3b;
  15'h7f28 : ret = 8'h10;
  15'h7f29 : ret = 8'h7b;
  15'h7f2a : ret = 8'hac;
  15'h7f2b : ret = 8'h3b;
  15'h7f2c : ret = 8'h11;
  15'h7f2d : ret = 8'h7b;
  15'h7f2e : ret = 8'hac;
  15'h7f2f : ret = 8'h3b;
  15'h7f30 : ret = 8'h18;
  15'h7f31 : ret = 8'h7b;
  15'h7f32 : ret = 8'h3d;
  15'h7f33 : ret = 8'h14;
  15'h7f34 : ret = 8'h3c;
  15'h7f35 : ret = 8'h10;
  15'h7f36 : ret = 8'h3b;
  15'h7f37 : ret = 8'h17;
  15'h7f38 : ret = 8'h7b;
  15'h7f39 : ret = 8'hac;
  15'h7f3a : ret = 8'h3b;
  15'h7f3b : ret = 8'h1f;
  15'h7f3c : ret = 8'h7b;
  15'h7f3d : ret = 8'hac;
  15'h7f3e : ret = 8'h3b;
  15'h7f3f : ret = 8'h14;
  15'h7f40 : ret = 8'h7b;
  15'h7f41 : ret = 8'hac;
  15'h7f42 : ret = 8'h3b;
  15'h7f43 : ret = 8'h16;
  15'h7f44 : ret = 8'h7b;
  15'h7f45 : ret = 8'h3a;
  15'h7f46 : ret = 8'h0;
  15'h7f47 : ret = 8'h10;
  15'h7f48 : ret = 8'hc1;
  15'h7f49 : ret = 8'h28;
  15'h7f4a : ret = 8'h9;
  15'h7f4b : ret = 8'h2a;
  15'h7f4c : ret = 8'h8;
  15'h7f4d : ret = 8'h11;
  15'h7f4e : ret = 8'h3d;
  15'h7f4f : ret = 8'h14;
  15'h7f50 : ret = 8'h3c;
  15'h7f51 : ret = 8'h10;
  15'h7f52 : ret = 8'h3b;
  15'h7f53 : ret = 8'h1f;
  15'h7f54 : ret = 8'h7b;
  15'h7f55 : ret = 8'hac;
  15'h7f56 : ret = 8'h3b;
  15'h7f57 : ret = 8'h1f;
  15'h7f58 : ret = 8'h7b;
  15'h7f59 : ret = 8'hac;
  15'h7f5a : ret = 8'h3b;
  15'h7f5b : ret = 8'h10;
  15'h7f5c : ret = 8'h7b;
  15'h7f5d : ret = 8'hac;
  15'h7f5e : ret = 8'h3b;
  15'h7f5f : ret = 8'h14;
  15'h7f60 : ret = 8'h7b;
  15'h7f61 : ret = 8'h31;
  15'h7f62 : ret = 8'h10;
  15'h7f63 : ret = 8'he1;
  15'h7f64 : ret = 8'h11;
  15'h7f65 : ret = 8'h41;
  15'h7f66 : ret = 8'h31;
  15'h7f67 : ret = 8'h10;
  15'h7f68 : ret = 8'he1;
  15'h7f69 : ret = 8'h11;
  15'h7f6a : ret = 8'h41;
  15'h7f6b : ret = 8'h31;
  15'h7f6c : ret = 8'h10;
  15'h7f6d : ret = 8'he1;
  15'h7f6e : ret = 8'h19;
  15'h7f6f : ret = 8'h41;
  15'h7f70 : ret = 8'h31;
  15'h7f71 : ret = 8'h10;
  15'h7f72 : ret = 8'he1;
  15'h7f73 : ret = 8'h11;
  15'h7f74 : ret = 8'h41;
  15'h7f75 : ret = 8'h31;
  15'h7f76 : ret = 8'h10;
  15'h7f77 : ret = 8'he1;
  15'h7f78 : ret = 8'h11;
  15'h7f79 : ret = 8'h41;
  15'h7f7a : ret = 8'h31;
  15'h7f7b : ret = 8'h10;
  15'h7f7c : ret = 8'he1;
  15'h7f7d : ret = 8'h11;
  15'h7f7e : ret = 8'h41;
  15'h7f7f : ret = 8'h31;
  15'h7f80 : ret = 8'h10;
  15'h7f81 : ret = 8'he1;
  15'h7f82 : ret = 8'h11;
  15'h7f83 : ret = 8'h41;
  15'h7f84 : ret = 8'h31;
  15'h7f85 : ret = 8'h10;
  15'h7f86 : ret = 8'he1;
  15'h7f87 : ret = 8'h11;
  15'h7f88 : ret = 8'h41;
  15'h7f89 : ret = 8'h31;
  15'h7f8a : ret = 8'h10;
  15'h7f8b : ret = 8'he1;
  15'h7f8c : ret = 8'h31;
  15'h7f8d : ret = 8'h32;
  15'h7f8e : ret = 8'h33;
  15'h7f8f : ret = 8'h34;
  15'h7f90 : ret = 8'h35;
  15'h7f91 : ret = 8'h36;
  15'h7f92 : ret = 8'h37;
  15'h7f93 : ret = 8'h38;
  15'h7f94 : ret = 8'h39;
  15'h7f95 : ret = 8'h3a;
  15'h7f96 : ret = 8'h3b;
  15'h7f97 : ret = 8'h3c;
  15'h7f98 : ret = 8'h3f;
  15'h7f99 : ret = 8'h14;
  15'h7f9a : ret = 8'h8;
  15'h7f9b : ret = 8'h34;
  15'h7f9c : ret = 8'h26;
  15'h7f9d : ret = 8'h31;
  15'h7f9e : ret = 8'h10;
  15'h7f9f : ret = 8'he3;
  15'h7fa0 : ret = 8'hf7;
  15'h7fa1 : ret = 8'he2;
  15'h7fa2 : ret = 8'h11;
  15'h7fa3 : ret = 8'h42;
  15'h7fa4 : ret = 8'h32;
  15'h7fa5 : ret = 8'h24;
  15'h7fa6 : ret = 8'h2;
  15'h7fa7 : ret = 8'h35;
  15'h7fa8 : ret = 8'h10;
  15'h7fa9 : ret = 8'he3;
  15'h7faa : ret = 8'h11;
  15'h7fab : ret = 8'h39;
  15'h7fac : ret = 8'h21;
  15'h7fad : ret = 8'h59;
  15'h7fae : ret = 8'h31;
  15'h7faf : ret = 8'h25;
  15'h7fb0 : ret = 8'h2;
  15'h7fb1 : ret = 8'h0;
  default: ret = 0;
endcase
endmodule
