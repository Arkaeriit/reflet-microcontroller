module rom10(input clk, input enable, input [14-1:0] addr, output [16-1:0] data);
    reg [16-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            14'h0 : data_reg <= 16'h5341;
            14'h1 : data_reg <= 16'h4D52;
            14'h2 : data_reg <= 16'h2D3C;
            14'h3 : data_reg <= 16'h2C3B;
            14'h4 : data_reg <= 16'h3D10;
            14'h5 : data_reg <= 16'h3C12;
            14'h6 : data_reg <= 16'h4C12;
            14'h7 : data_reg <= 16'h3E4E;
            14'h8 : data_reg <= 16'h8000;
            14'h9 : data_reg <= 16'h4C13;
            14'hA : data_reg <= 16'h4E08;
            14'hB : data_reg <= 16'h3CF0;
            14'hC : data_reg <= 16'h3D2B;
            14'hD : data_reg <= 16'h3F2C;
            14'hE : data_reg <= 16'h2D3C;
            14'hF : data_reg <= 16'h2C3B;
            14'h10 : data_reg <= 16'h3D10;
            14'h11 : data_reg <= 16'h3C12;
            14'h12 : data_reg <= 16'h4C12;
            14'h13 : data_reg <= 16'h3E4E;
            14'h14 : data_reg <= 16'h023D;
            14'h15 : data_reg <= 16'h4C13;
            14'h16 : data_reg <= 16'h4E08;
            14'h17 : data_reg <= 16'h3CF0;
            14'h18 : data_reg <= 16'h3D2B;
            14'h19 : data_reg <= 16'h3E2C;
            14'h1A : data_reg <= 16'h233C;
            14'h1B : data_reg <= 16'h2C0B;
            14'h1C : data_reg <= 16'h243C;
            14'h1D : data_reg <= 16'h2C0B;
            14'h1E : data_reg <= 16'h253C;
            14'h1F : data_reg <= 16'h2C0B;
            14'h20 : data_reg <= 16'h263C;
            14'h21 : data_reg <= 16'h2C0B;
            14'h22 : data_reg <= 16'h3310;
            14'h23 : data_reg <= 16'h3C34;
            14'h24 : data_reg <= 16'h3B2D;
            14'h25 : data_reg <= 16'h102C;
            14'h26 : data_reg <= 16'h123D;
            14'h27 : data_reg <= 16'h003C;
            14'h28 : data_reg <= 16'h4C12;
            14'h29 : data_reg <= 16'h3E4E;
            14'h2A : data_reg <= 16'h0085;
            14'h2B : data_reg <= 16'h4C13;
            14'h2C : data_reg <= 16'h4E08;
            14'h2D : data_reg <= 16'h3CF0;
            14'h2E : data_reg <= 16'h3D2B;
            14'h2F : data_reg <= 16'h352C;
            14'h30 : data_reg <= 16'h2D3C;
            14'h31 : data_reg <= 16'h2C3B;
            14'h32 : data_reg <= 16'h3D10;
            14'h33 : data_reg <= 16'h3C12;
            14'h34 : data_reg <= 16'h4C12;
            14'h35 : data_reg <= 16'h3E4E;
            14'h36 : data_reg <= 16'h0079;
            14'h37 : data_reg <= 16'h4C13;
            14'h38 : data_reg <= 16'h4E08;
            14'h39 : data_reg <= 16'h3CF0;
            14'h3A : data_reg <= 16'h3D2B;
            14'h3B : data_reg <= 16'h362C;
            14'h3C : data_reg <= 16'h2410;
            14'h3D : data_reg <= 16'h25C2;
            14'h3E : data_reg <= 16'h1109;
            14'h3F : data_reg <= 16'h3444;
            14'h40 : data_reg <= 16'h4321;
            14'h41 : data_reg <= 16'h2633;
            14'h42 : data_reg <= 16'h233E;
            14'h43 : data_reg <= 16'h3C31;
            14'h44 : data_reg <= 16'h360A;
            14'h45 : data_reg <= 16'h3C2C;
            14'h46 : data_reg <= 16'h350A;
            14'h47 : data_reg <= 16'h3C2C;
            14'h48 : data_reg <= 16'h340A;
            14'h49 : data_reg <= 16'h3C2C;
            14'h4A : data_reg <= 16'h330A;
            14'h4B : data_reg <= 16'h0D2C;
            14'h4C : data_reg <= 16'h233C;
            14'h4D : data_reg <= 16'h2C0B;
            14'h4E : data_reg <= 16'h253C;
            14'h4F : data_reg <= 16'h2C0B;
            14'h50 : data_reg <= 16'h263C;
            14'h51 : data_reg <= 16'h2C0B;
            14'h52 : data_reg <= 16'h2D3C;
            14'h53 : data_reg <= 16'h2C3B;
            14'h54 : data_reg <= 16'h3D10;
            14'h55 : data_reg <= 16'h3C12;
            14'h56 : data_reg <= 16'h4C12;
            14'h57 : data_reg <= 16'h3E4E;
            14'h58 : data_reg <= 16'h00D6;
            14'h59 : data_reg <= 16'h4C13;
            14'h5A : data_reg <= 16'h4E08;
            14'h5B : data_reg <= 16'h3CF0;
            14'h5C : data_reg <= 16'h3D2B;
            14'h5D : data_reg <= 16'h352C;
            14'h5E : data_reg <= 16'h2D3C;
            14'h5F : data_reg <= 16'h2C3B;
            14'h60 : data_reg <= 16'h3D10;
            14'h61 : data_reg <= 16'h3C12;
            14'h62 : data_reg <= 16'h4C12;
            14'h63 : data_reg <= 16'h3E4E;
            14'h64 : data_reg <= 16'h00E2;
            14'h65 : data_reg <= 16'h4C13;
            14'h66 : data_reg <= 16'h4E08;
            14'h67 : data_reg <= 16'h3CF0;
            14'h68 : data_reg <= 16'h3D2B;
            14'h69 : data_reg <= 16'h362C;
            14'h6A : data_reg <= 16'h3310;
            14'h6B : data_reg <= 16'hD221;
            14'h6C : data_reg <= 16'h0926;
            14'h6D : data_reg <= 16'h5221;
            14'h6E : data_reg <= 16'h1131;
            14'h6F : data_reg <= 16'h3343;
            14'h70 : data_reg <= 16'h3E25;
            14'h71 : data_reg <= 16'h3221;
            14'h72 : data_reg <= 16'h3123;
            14'h73 : data_reg <= 16'h0A3C;
            14'h74 : data_reg <= 16'h2C36;
            14'h75 : data_reg <= 16'h0A3C;
            14'h76 : data_reg <= 16'h2C35;
            14'h77 : data_reg <= 16'h0A3C;
            14'h78 : data_reg <= 16'h2C33;
            14'h79 : data_reg <= 16'h3C0D;
            14'h7A : data_reg <= 16'h0B23;
            14'h7B : data_reg <= 16'h3C2C;
            14'h7C : data_reg <= 16'h0B24;
            14'h7D : data_reg <= 16'h3C2C;
            14'h7E : data_reg <= 16'h0B25;
            14'h7F : data_reg <= 16'h3C2C;
            14'h80 : data_reg <= 16'h0B26;
            14'h81 : data_reg <= 16'h3C2C;
            14'h82 : data_reg <= 16'h0B27;
            14'h83 : data_reg <= 16'h3C2C;
            14'h84 : data_reg <= 16'h3B2D;
            14'h85 : data_reg <= 16'h102C;
            14'h86 : data_reg <= 16'h123D;
            14'h87 : data_reg <= 16'h003C;
            14'h88 : data_reg <= 16'h4C12;
            14'h89 : data_reg <= 16'h3E4E;
            14'h8A : data_reg <= 16'h0173;
            14'h8B : data_reg <= 16'h4C13;
            14'h8C : data_reg <= 16'h4E08;
            14'h8D : data_reg <= 16'h3CF0;
            14'h8E : data_reg <= 16'h3D2B;
            14'h8F : data_reg <= 16'h352C;
            14'h90 : data_reg <= 16'h2D3C;
            14'h91 : data_reg <= 16'h2C3B;
            14'h92 : data_reg <= 16'h3D10;
            14'h93 : data_reg <= 16'h3C12;
            14'h94 : data_reg <= 16'h4C12;
            14'h95 : data_reg <= 16'h3E4E;
            14'h96 : data_reg <= 16'h0154;
            14'h97 : data_reg <= 16'h4C13;
            14'h98 : data_reg <= 16'h4E08;
            14'h99 : data_reg <= 16'h3CF0;
            14'h9A : data_reg <= 16'h3D2B;
            14'h9B : data_reg <= 16'h362C;
            14'h9C : data_reg <= 16'h2D3C;
            14'h9D : data_reg <= 16'h2C3B;
            14'h9E : data_reg <= 16'h3D10;
            14'h9F : data_reg <= 16'h3C12;
            14'hA0 : data_reg <= 16'h4C12;
            14'hA1 : data_reg <= 16'h3E4E;
            14'hA2 : data_reg <= 16'h0034;
            14'hA3 : data_reg <= 16'h4C13;
            14'hA4 : data_reg <= 16'h4E08;
            14'hA5 : data_reg <= 16'h3CF0;
            14'hA6 : data_reg <= 16'h3D2B;
            14'hA7 : data_reg <= 16'h372C;
            14'hA8 : data_reg <= 16'h3311;
            14'hA9 : data_reg <= 16'h3410;
            14'hAA : data_reg <= 16'hC224;
            14'hAB : data_reg <= 16'h0925;
            14'hAC : data_reg <= 16'h4411;
            14'hAD : data_reg <= 16'h3C34;
            14'hAE : data_reg <= 16'h0B21;
            14'hAF : data_reg <= 16'h3C2C;
            14'hB0 : data_reg <= 16'h0B22;
            14'hB1 : data_reg <= 16'h232C;
            14'hB2 : data_reg <= 16'h2732;
            14'hB3 : data_reg <= 16'h210C;
            14'hB4 : data_reg <= 16'h3C33;
            14'hB5 : data_reg <= 16'h320A;
            14'hB6 : data_reg <= 16'h3C2C;
            14'hB7 : data_reg <= 16'h310A;
            14'hB8 : data_reg <= 16'h262C;
            14'hB9 : data_reg <= 16'h233E;
            14'hBA : data_reg <= 16'h3C31;
            14'hBB : data_reg <= 16'h370A;
            14'hBC : data_reg <= 16'h3C2C;
            14'hBD : data_reg <= 16'h360A;
            14'hBE : data_reg <= 16'h3C2C;
            14'hBF : data_reg <= 16'h350A;
            14'hC0 : data_reg <= 16'h3C2C;
            14'hC1 : data_reg <= 16'h340A;
            14'hC2 : data_reg <= 16'h3C2C;
            14'hC3 : data_reg <= 16'h330A;
            14'hC4 : data_reg <= 16'h0D2C;
            14'hC5 : data_reg <= 16'h7D00;
            14'hC6 : data_reg <= 16'h8000;
            14'hC7 : data_reg <= 16'hFF00;
            14'hC8 : data_reg <= 16'hFF04;
            14'hC9 : data_reg <= 16'hFF08;
            14'hCA : data_reg <= 16'hFF10;
            14'hCB : data_reg <= 16'hFF13;
            14'hCC : data_reg <= 16'hFF16;
            14'hCD : data_reg <= 16'hFF1A;
            14'hCE : data_reg <= 16'hFF1C;
            14'hCF : data_reg <= 16'hFF1F;
            14'hD0 : data_reg <= 16'hFF21;
            14'hD1 : data_reg <= 16'hFF22;
            14'hD2 : data_reg <= 16'h4121;
            14'hD3 : data_reg <= 16'h314A;
            14'hD4 : data_reg <= 16'h210D;
            14'hD5 : data_reg <= 16'h110B;
            14'hD6 : data_reg <= 16'hFA31;
            14'hD7 : data_reg <= 16'h0C0F;
            14'hD8 : data_reg <= 16'h31F1;
            14'hD9 : data_reg <= 16'h2D0F;
            14'hDA : data_reg <= 16'h160B;
            14'hDB : data_reg <= 16'h223D;
            14'hDC : data_reg <= 16'h11E1;
            14'hDD : data_reg <= 16'h3141;
            14'hDE : data_reg <= 16'h2331;
            14'hDF : data_reg <= 16'h11E1;
            14'hE0 : data_reg <= 16'h3141;
            14'hE1 : data_reg <= 16'h2431;
            14'hE2 : data_reg <= 16'h0AE1;
            14'hE3 : data_reg <= 16'h0A3D;
            14'hE4 : data_reg <= 16'h0D31;
            14'hE5 : data_reg <= 16'h0B21;
            14'hE6 : data_reg <= 16'h312A;
            14'hE7 : data_reg <= 16'h3C0F;
            14'hE8 : data_reg <= 16'h3B2D;
            14'hE9 : data_reg <= 16'h102C;
            14'hEA : data_reg <= 16'h123D;
            14'hEB : data_reg <= 16'h003C;
            14'hEC : data_reg <= 16'h4C12;
            14'hED : data_reg <= 16'h3E4E;
            14'hEE : data_reg <= 16'h01A4;
            14'hEF : data_reg <= 16'h4C13;
            14'hF0 : data_reg <= 16'h4E08;
            14'hF1 : data_reg <= 16'h3CF0;
            14'hF2 : data_reg <= 16'h3D2B;
            14'hF3 : data_reg <= 16'hE12C;
            14'hF4 : data_reg <= 16'h4112;
            14'hF5 : data_reg <= 16'h0F31;
            14'hF6 : data_reg <= 16'h2D3C;
            14'hF7 : data_reg <= 16'h2C3B;
            14'hF8 : data_reg <= 16'h3D10;
            14'hF9 : data_reg <= 16'h3C12;
            14'hFA : data_reg <= 16'h4C12;
            14'hFB : data_reg <= 16'h3E4E;
            14'hFC : data_reg <= 16'hFF24;
            14'hFD : data_reg <= 16'h4C13;
            14'hFE : data_reg <= 16'h4E08;
            14'hFF : data_reg <= 16'h3CF0;
            14'h100 : data_reg <= 16'h3D2B;
            14'h101 : data_reg <= 16'hE12C;
            14'h102 : data_reg <= 16'h4112;
            14'h103 : data_reg <= 16'h0F31;
            14'h104 : data_reg <= 16'h2D3C;
            14'h105 : data_reg <= 16'h2C3B;
            14'h106 : data_reg <= 16'h3D10;
            14'h107 : data_reg <= 16'h3C12;
            14'h108 : data_reg <= 16'h4C12;
            14'h109 : data_reg <= 16'h3E4E;
            14'h10A : data_reg <= 16'h01A9;
            14'h10B : data_reg <= 16'h4C13;
            14'h10C : data_reg <= 16'h4E08;
            14'h10D : data_reg <= 16'h3CF0;
            14'h10E : data_reg <= 16'h3D2B;
            14'h10F : data_reg <= 16'hE12C;
            14'h110 : data_reg <= 16'h4112;
            14'h111 : data_reg <= 16'h0F31;
            14'h112 : data_reg <= 16'h3C14;
            14'h113 : data_reg <= 16'hAC1A;
            14'h114 : data_reg <= 16'h103C;
            14'h115 : data_reg <= 16'hE17C;
            14'h116 : data_reg <= 16'h4112;
            14'h117 : data_reg <= 16'h0F31;
            14'h118 : data_reg <= 16'h3C14;
            14'h119 : data_reg <= 16'hAC17;
            14'h11A : data_reg <= 16'h183C;
            14'h11B : data_reg <= 16'hE17C;
            14'h11C : data_reg <= 16'h0A3C;
            14'h11D : data_reg <= 16'h2C31;
            14'h11E : data_reg <= 16'h120D;
            14'h11F : data_reg <= 16'h1531;
            14'h120 : data_reg <= 16'h3C32;
            14'h121 : data_reg <= 16'h3B2D;
            14'h122 : data_reg <= 16'h102C;
            14'h123 : data_reg <= 16'h123D;
            14'h124 : data_reg <= 16'h003C;
            14'h125 : data_reg <= 16'h4C12;
            14'h126 : data_reg <= 16'h3E4E;
            14'h127 : data_reg <= 16'h0034;
            14'h128 : data_reg <= 16'h4C13;
            14'h129 : data_reg <= 16'h4E08;
            14'h12A : data_reg <= 16'h3CF0;
            14'h12B : data_reg <= 16'h3D2B;
            14'h12C : data_reg <= 16'h0C2C;
            14'h12D : data_reg <= 16'h3A2F;
            14'h12E : data_reg <= 16'h3F41;
            14'h12F : data_reg <= 16'h2D3C;
            14'h130 : data_reg <= 16'h2C3B;
            14'h131 : data_reg <= 16'h3D10;
            14'h132 : data_reg <= 16'h3C12;
            14'h133 : data_reg <= 16'h4C12;
            14'h134 : data_reg <= 16'h3E4E;
            14'h135 : data_reg <= 16'h01CA;
            14'h136 : data_reg <= 16'h4C13;
            14'h137 : data_reg <= 16'h4E08;
            14'h138 : data_reg <= 16'h3CF0;
            14'h139 : data_reg <= 16'h3D2B;
            14'h13A : data_reg <= 16'h0C2C;
            14'h13B : data_reg <= 16'h3C14;
            14'h13C : data_reg <= 16'hAC10;
            14'h13D : data_reg <= 16'h1A3C;
            14'h13E : data_reg <= 16'h327C;
            14'h13F : data_reg <= 16'h3C14;
            14'h140 : data_reg <= 16'hAC10;
            14'h141 : data_reg <= 16'h1A3C;
            14'h142 : data_reg <= 16'h337C;
            14'h143 : data_reg <= 16'h3413;
            14'h144 : data_reg <= 16'h2D3C;
            14'h145 : data_reg <= 16'h2C3B;
            14'h146 : data_reg <= 16'h3D10;
            14'h147 : data_reg <= 16'h3C12;
            14'h148 : data_reg <= 16'h4C12;
            14'h149 : data_reg <= 16'h3E4E;
            14'h14A : data_reg <= 16'h01A9;
            14'h14B : data_reg <= 16'h4C13;
            14'h14C : data_reg <= 16'h4E08;
            14'h14D : data_reg <= 16'h3CF0;
            14'h14E : data_reg <= 16'h3D2B;
            14'h14F : data_reg <= 16'h0C2C;
            14'h150 : data_reg <= 16'h113C;
            14'h151 : data_reg <= 16'h3242;
            14'h152 : data_reg <= 16'h2C32;
            14'h153 : data_reg <= 16'h2D3C;
            14'h154 : data_reg <= 16'h2C3B;
            14'h155 : data_reg <= 16'h3D10;
            14'h156 : data_reg <= 16'h3C12;
            14'h157 : data_reg <= 16'h4C12;
            14'h158 : data_reg <= 16'h3E4E;
            14'h159 : data_reg <= 16'h01A9;
            14'h15A : data_reg <= 16'h4C13;
            14'h15B : data_reg <= 16'h4E08;
            14'h15C : data_reg <= 16'h3CF0;
            14'h15D : data_reg <= 16'h3D2B;
            14'h15E : data_reg <= 16'h0C2C;
            14'h15F : data_reg <= 16'h113C;
            14'h160 : data_reg <= 16'h3242;
            14'h161 : data_reg <= 16'h2C32;
            14'h162 : data_reg <= 16'h2D3C;
            14'h163 : data_reg <= 16'h2C3B;
            14'h164 : data_reg <= 16'h3D10;
            14'h165 : data_reg <= 16'h3C12;
            14'h166 : data_reg <= 16'h4C12;
            14'h167 : data_reg <= 16'h3E4E;
            14'h168 : data_reg <= 16'h01A9;
            14'h169 : data_reg <= 16'h4C13;
            14'h16A : data_reg <= 16'h4E08;
            14'h16B : data_reg <= 16'h3CF0;
            14'h16C : data_reg <= 16'h3D2B;
            14'h16D : data_reg <= 16'h0C2C;
            14'h16E : data_reg <= 16'h113C;
            14'h16F : data_reg <= 16'h3242;
            14'h170 : data_reg <= 16'h2C32;
            14'h171 : data_reg <= 16'h2D3C;
            14'h172 : data_reg <= 16'h2C3B;
            14'h173 : data_reg <= 16'h3D10;
            14'h174 : data_reg <= 16'h3C12;
            14'h175 : data_reg <= 16'h4C12;
            14'h176 : data_reg <= 16'h3E4E;
            14'h177 : data_reg <= 16'h01A9;
            14'h178 : data_reg <= 16'h4C13;
            14'h179 : data_reg <= 16'h4E08;
            14'h17A : data_reg <= 16'h3CF0;
            14'h17B : data_reg <= 16'h3D2B;
            14'h17C : data_reg <= 16'h0C2C;
            14'h17D : data_reg <= 16'h113C;
            14'h17E : data_reg <= 16'h3242;
            14'h17F : data_reg <= 16'h2C32;
            14'h180 : data_reg <= 16'h2D3C;
            14'h181 : data_reg <= 16'h2C3B;
            14'h182 : data_reg <= 16'h3D10;
            14'h183 : data_reg <= 16'h3C12;
            14'h184 : data_reg <= 16'h4C12;
            14'h185 : data_reg <= 16'h3E4E;
            14'h186 : data_reg <= 16'h01A9;
            14'h187 : data_reg <= 16'h4C13;
            14'h188 : data_reg <= 16'h4E08;
            14'h189 : data_reg <= 16'h3CF0;
            14'h18A : data_reg <= 16'h3D2B;
            14'h18B : data_reg <= 16'h0C2C;
            14'h18C : data_reg <= 16'h113C;
            14'h18D : data_reg <= 16'h3242;
            14'h18E : data_reg <= 16'h2C32;
            14'h18F : data_reg <= 16'h2D3C;
            14'h190 : data_reg <= 16'h2C3B;
            14'h191 : data_reg <= 16'h3D10;
            14'h192 : data_reg <= 16'h3C12;
            14'h193 : data_reg <= 16'h4C12;
            14'h194 : data_reg <= 16'h3E4E;
            14'h195 : data_reg <= 16'h01A9;
            14'h196 : data_reg <= 16'h4C13;
            14'h197 : data_reg <= 16'h4E08;
            14'h198 : data_reg <= 16'h3CF0;
            14'h199 : data_reg <= 16'h3D2B;
            14'h19A : data_reg <= 16'h0C2C;
            14'h19B : data_reg <= 16'h113C;
            14'h19C : data_reg <= 16'h3242;
            14'h19D : data_reg <= 16'h2C32;
            14'h19E : data_reg <= 16'h2D3C;
            14'h19F : data_reg <= 16'h2C3B;
            14'h1A0 : data_reg <= 16'h3D10;
            14'h1A1 : data_reg <= 16'h3C12;
            14'h1A2 : data_reg <= 16'h4C12;
            14'h1A3 : data_reg <= 16'h3E4E;
            14'h1A4 : data_reg <= 16'h01A9;
            14'h1A5 : data_reg <= 16'h4C13;
            14'h1A6 : data_reg <= 16'h4E08;
            14'h1A7 : data_reg <= 16'h3CF0;
            14'h1A8 : data_reg <= 16'h3D2B;
            14'h1A9 : data_reg <= 16'h0C2C;
            14'h1AA : data_reg <= 16'h000E;
            default : data_reg <= 0;
        endcase
    assign data = ( enable ? data_reg : 0 );
endmodule
