../cpu/reflet.vh