module rom02(input clk, input enable, input [14-1:0] addr, output [16-1:0] data);
    reg [16-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            14'h0 : data_reg <= 16'h5341;
            14'h1 : data_reg <= 16'h4D52;
            14'h2 : data_reg <= 16'h2D3C;
            14'h3 : data_reg <= 16'h2C3B;
            14'h4 : data_reg <= 16'h3D10;
            14'h5 : data_reg <= 16'h3C12;
            14'h6 : data_reg <= 16'h4C12;
            14'h7 : data_reg <= 16'h3E4E;
            14'h8 : data_reg <= 16'h8000;
            14'h9 : data_reg <= 16'h4C13;
            14'hA : data_reg <= 16'h4E08;
            14'hB : data_reg <= 16'h3CF0;
            14'hC : data_reg <= 16'h3D2B;
            14'hD : data_reg <= 16'h3F2C;
            14'hE : data_reg <= 16'h2D3C;
            14'hF : data_reg <= 16'h2C3B;
            14'h10 : data_reg <= 16'h3D10;
            14'h11 : data_reg <= 16'h3C12;
            14'h12 : data_reg <= 16'h4C12;
            14'h13 : data_reg <= 16'h3E4E;
            14'h14 : data_reg <= 16'h0674;
            14'h15 : data_reg <= 16'h4C13;
            14'h16 : data_reg <= 16'h4E08;
            14'h17 : data_reg <= 16'h3CF0;
            14'h18 : data_reg <= 16'h3D2B;
            14'h19 : data_reg <= 16'h3E2C;
            14'h1A : data_reg <= 16'h223C;
            14'h1B : data_reg <= 16'h2C0B;
            14'h1C : data_reg <= 16'h243C;
            14'h1D : data_reg <= 16'h2C0B;
            14'h1E : data_reg <= 16'h2D3C;
            14'h1F : data_reg <= 16'h2C3B;
            14'h20 : data_reg <= 16'h3D10;
            14'h21 : data_reg <= 16'h3C12;
            14'h22 : data_reg <= 16'h4C12;
            14'h23 : data_reg <= 16'h3E4E;
            14'h24 : data_reg <= 16'h012A;
            14'h25 : data_reg <= 16'h4C13;
            14'h26 : data_reg <= 16'h4E08;
            14'h27 : data_reg <= 16'h3CF0;
            14'h28 : data_reg <= 16'h3D2B;
            14'h29 : data_reg <= 16'hF02C;
            14'h2A : data_reg <= 16'h3203;
            14'h2B : data_reg <= 16'h2D3C;
            14'h2C : data_reg <= 16'h2C3B;
            14'h2D : data_reg <= 16'h3D10;
            14'h2E : data_reg <= 16'h3C12;
            14'h2F : data_reg <= 16'h4C12;
            14'h30 : data_reg <= 16'h3E4E;
            14'h31 : data_reg <= 16'h006E;
            14'h32 : data_reg <= 16'h4C13;
            14'h33 : data_reg <= 16'h4E08;
            14'h34 : data_reg <= 16'h3CF0;
            14'h35 : data_reg <= 16'h3D2B;
            14'h36 : data_reg <= 16'h342C;
            14'h37 : data_reg <= 16'h3CF2;
            14'h38 : data_reg <= 16'hCC10;
            14'h39 : data_reg <= 16'h0924;
            14'h3A : data_reg <= 16'h4211;
            14'h3B : data_reg <= 16'h213C;
            14'h3C : data_reg <= 16'h10EC;
            14'h3D : data_reg <= 16'h03E2;
            14'h3E : data_reg <= 16'h0A3C;
            14'h3F : data_reg <= 16'h2C34;
            14'h40 : data_reg <= 16'h0A3C;
            14'h41 : data_reg <= 16'h2C32;
            14'h42 : data_reg <= 16'h3C0D;
            14'h43 : data_reg <= 16'h0B21;
            14'h44 : data_reg <= 16'h1A2C;
            14'h45 : data_reg <= 16'h3C31;
            14'h46 : data_reg <= 16'h3B2D;
            14'h47 : data_reg <= 16'h102C;
            14'h48 : data_reg <= 16'h123D;
            14'h49 : data_reg <= 16'h003C;
            14'h4A : data_reg <= 16'h4C12;
            14'h4B : data_reg <= 16'h3E4E;
            14'h4C : data_reg <= 16'h0034;
            14'h4D : data_reg <= 16'h4C13;
            14'h4E : data_reg <= 16'h4E08;
            14'h4F : data_reg <= 16'h3CF0;
            14'h50 : data_reg <= 16'h3D2B;
            14'h51 : data_reg <= 16'h0C2C;
            14'h52 : data_reg <= 16'h311D;
            14'h53 : data_reg <= 16'h2D3C;
            14'h54 : data_reg <= 16'h2C3B;
            14'h55 : data_reg <= 16'h3D10;
            14'h56 : data_reg <= 16'h3C12;
            14'h57 : data_reg <= 16'h4C12;
            14'h58 : data_reg <= 16'h3E4E;
            14'h59 : data_reg <= 16'h0034;
            14'h5A : data_reg <= 16'h4C13;
            14'h5B : data_reg <= 16'h4E08;
            14'h5C : data_reg <= 16'h3CF0;
            14'h5D : data_reg <= 16'h3D2B;
            14'h5E : data_reg <= 16'h0C2C;
            14'h5F : data_reg <= 16'h0A3C;
            14'h60 : data_reg <= 16'h2C31;
            14'h61 : data_reg <= 16'h3C0D;
            14'h62 : data_reg <= 16'h0B22;
            14'h63 : data_reg <= 16'h3C2C;
            14'h64 : data_reg <= 16'h0B23;
            14'h65 : data_reg <= 16'h3C2C;
            14'h66 : data_reg <= 16'h3B2D;
            14'h67 : data_reg <= 16'h102C;
            14'h68 : data_reg <= 16'h123D;
            14'h69 : data_reg <= 16'h003C;
            14'h6A : data_reg <= 16'h4C12;
            14'h6B : data_reg <= 16'h3E4E;
            14'h6C : data_reg <= 16'h012A;
            14'h6D : data_reg <= 16'h4C13;
            14'h6E : data_reg <= 16'h4E08;
            14'h6F : data_reg <= 16'h3CF0;
            14'h70 : data_reg <= 16'h3D2B;
            14'h71 : data_reg <= 16'hF02C;
            14'h72 : data_reg <= 16'h1232;
            14'h73 : data_reg <= 16'h3242;
            14'h74 : data_reg <= 16'h2D3C;
            14'h75 : data_reg <= 16'h2C3B;
            14'h76 : data_reg <= 16'h3D10;
            14'h77 : data_reg <= 16'h3C12;
            14'h78 : data_reg <= 16'h4C12;
            14'h79 : data_reg <= 16'h3E4E;
            14'h7A : data_reg <= 16'h0105;
            14'h7B : data_reg <= 16'h4C13;
            14'h7C : data_reg <= 16'h4E08;
            14'h7D : data_reg <= 16'h3CF0;
            14'h7E : data_reg <= 16'h3D2B;
            14'h7F : data_reg <= 16'h332C;
            14'h80 : data_reg <= 16'h0311;
            14'h81 : data_reg <= 16'h03E2;
            14'h82 : data_reg <= 16'h0331;
            14'h83 : data_reg <= 16'h03F2;
            14'h84 : data_reg <= 16'h23C1;
            14'h85 : data_reg <= 16'h1109;
            14'h86 : data_reg <= 16'h3242;
            14'h87 : data_reg <= 16'hF203;
            14'h88 : data_reg <= 16'h3103;
            14'h89 : data_reg <= 16'h0A3C;
            14'h8A : data_reg <= 16'h2C33;
            14'h8B : data_reg <= 16'h0A3C;
            14'h8C : data_reg <= 16'h2C32;
            14'h8D : data_reg <= 16'h000D;
            14'h8E : data_reg <= 16'h7D00;
            14'h8F : data_reg <= 16'h8000;
            14'h90 : data_reg <= 16'hFF00;
            14'h91 : data_reg <= 16'hFF04;
            14'h92 : data_reg <= 16'hFF08;
            14'h93 : data_reg <= 16'hFF10;
            14'h94 : data_reg <= 16'hFF13;
            14'h95 : data_reg <= 16'hFF16;
            14'h96 : data_reg <= 16'hFF1A;
            14'h97 : data_reg <= 16'hFF1C;
            14'h98 : data_reg <= 16'hFF1F;
            14'h99 : data_reg <= 16'hFF21;
            14'h9A : data_reg <= 16'hFF22;
            14'h9B : data_reg <= 16'h213C;
            14'h9C : data_reg <= 16'h2C0B;
            14'h9D : data_reg <= 16'h223C;
            14'h9E : data_reg <= 16'h2C0B;
            14'h9F : data_reg <= 16'h233C;
            14'hA0 : data_reg <= 16'h2C0B;
            14'hA1 : data_reg <= 16'h243C;
            14'hA2 : data_reg <= 16'h2C0B;
            14'hA3 : data_reg <= 16'h253C;
            14'hA4 : data_reg <= 16'h2C0B;
            14'hA5 : data_reg <= 16'h263C;
            14'hA6 : data_reg <= 16'h2C0B;
            14'hA7 : data_reg <= 16'h2D3C;
            14'hA8 : data_reg <= 16'h2C3B;
            14'hA9 : data_reg <= 16'h3D10;
            14'hAA : data_reg <= 16'h3C12;
            14'hAB : data_reg <= 16'h4C12;
            14'hAC : data_reg <= 16'h3E4E;
            14'hAD : data_reg <= 16'h0198;
            14'hAE : data_reg <= 16'h4C13;
            14'hAF : data_reg <= 16'h4E08;
            14'hB0 : data_reg <= 16'h3CF0;
            14'hB1 : data_reg <= 16'h3D2B;
            14'hB2 : data_reg <= 16'h332C;
            14'hB3 : data_reg <= 16'h2D3C;
            14'hB4 : data_reg <= 16'h2C3B;
            14'hB5 : data_reg <= 16'h3D10;
            14'hB6 : data_reg <= 16'h3C12;
            14'hB7 : data_reg <= 16'h4C12;
            14'hB8 : data_reg <= 16'h3E4E;
            14'hB9 : data_reg <= 16'h01B6;
            14'hBA : data_reg <= 16'h4C13;
            14'hBB : data_reg <= 16'h4E08;
            14'hBC : data_reg <= 16'h3CF0;
            14'hBD : data_reg <= 16'h3D2B;
            14'hBE : data_reg <= 16'h342C;
            14'hBF : data_reg <= 16'h3511;
            14'hC0 : data_reg <= 16'h2D3C;
            14'hC1 : data_reg <= 16'h2C3B;
            14'hC2 : data_reg <= 16'h3D10;
            14'hC3 : data_reg <= 16'h3C12;
            14'hC4 : data_reg <= 16'h4C12;
            14'hC5 : data_reg <= 16'h3E4E;
            14'hC6 : data_reg <= 16'h0034;
            14'hC7 : data_reg <= 16'h4C13;
            14'hC8 : data_reg <= 16'h4E08;
            14'hC9 : data_reg <= 16'h3CF0;
            14'hCA : data_reg <= 16'h3D2B;
            14'hCB : data_reg <= 16'h362C;
            14'hCC : data_reg <= 16'hC210;
            14'hCD : data_reg <= 16'h0924;
            14'hCE : data_reg <= 16'hF103;
            14'hCF : data_reg <= 16'h3C03;
            14'hD0 : data_reg <= 16'h213C;
            14'hD1 : data_reg <= 16'h2C0B;
            14'hD2 : data_reg <= 16'h2C3C;
            14'hD3 : data_reg <= 16'h2C31;
            14'hD4 : data_reg <= 16'h0C26;
            14'hD5 : data_reg <= 16'h0A3C;
            14'hD6 : data_reg <= 16'h2C31;
            14'hD7 : data_reg <= 16'h4521;
            14'hD8 : data_reg <= 16'h2231;
            14'hD9 : data_reg <= 16'h3255;
            14'hDA : data_reg <= 16'h3E23;
            14'hDB : data_reg <= 16'h0A3C;
            14'hDC : data_reg <= 16'h2C36;
            14'hDD : data_reg <= 16'h0A3C;
            14'hDE : data_reg <= 16'h2C35;
            14'hDF : data_reg <= 16'h0A3C;
            14'hE0 : data_reg <= 16'h2C34;
            14'hE1 : data_reg <= 16'h0A3C;
            14'hE2 : data_reg <= 16'h2C33;
            14'hE3 : data_reg <= 16'h0A3C;
            14'hE4 : data_reg <= 16'h2C32;
            14'hE5 : data_reg <= 16'h0A3C;
            14'hE6 : data_reg <= 16'h2C31;
            14'hE7 : data_reg <= 16'h3C0D;
            14'hE8 : data_reg <= 16'h0B22;
            14'hE9 : data_reg <= 16'h3C2C;
            14'hEA : data_reg <= 16'h0B21;
            14'hEB : data_reg <= 16'h3C2C;
            14'hEC : data_reg <= 16'h3B2D;
            14'hED : data_reg <= 16'h102C;
            14'hEE : data_reg <= 16'h123D;
            14'hEF : data_reg <= 16'h003C;
            14'hF0 : data_reg <= 16'h4C12;
            14'hF1 : data_reg <= 16'h3E4E;
            14'hF2 : data_reg <= 16'h04E2;
            14'hF3 : data_reg <= 16'h4C13;
            14'hF4 : data_reg <= 16'h4E08;
            14'hF5 : data_reg <= 16'h3CF0;
            14'hF6 : data_reg <= 16'h3D2B;
            14'hF7 : data_reg <= 16'h0C2C;
            14'hF8 : data_reg <= 16'h213C;
            14'hF9 : data_reg <= 16'h2C32;
            14'hFA : data_reg <= 16'h0A3C;
            14'hFB : data_reg <= 16'h2C31;
            14'hFC : data_reg <= 16'h2D3C;
            14'hFD : data_reg <= 16'h2C3B;
            14'hFE : data_reg <= 16'h3D10;
            14'hFF : data_reg <= 16'h3C12;
            14'h100 : data_reg <= 16'h4C12;
            14'h101 : data_reg <= 16'h3E4E;
            14'h102 : data_reg <= 16'h0136;
            14'h103 : data_reg <= 16'h4C13;
            14'h104 : data_reg <= 16'h4E08;
            14'h105 : data_reg <= 16'h3CF0;
            14'h106 : data_reg <= 16'h3D2B;
            14'h107 : data_reg <= 16'h0C2C;
            14'h108 : data_reg <= 16'h0A3C;
            14'h109 : data_reg <= 16'h2C32;
            14'h10A : data_reg <= 16'h100D;
            14'h10B : data_reg <= 16'h3CC1;
            14'h10C : data_reg <= 16'h3B2D;
            14'h10D : data_reg <= 16'h102C;
            14'h10E : data_reg <= 16'h123D;
            14'h10F : data_reg <= 16'h003C;
            14'h110 : data_reg <= 16'h4C12;
            14'h111 : data_reg <= 16'h3E4E;
            14'h112 : data_reg <= 16'h030F;
            14'h113 : data_reg <= 16'h4C13;
            14'h114 : data_reg <= 16'h4E08;
            14'h115 : data_reg <= 16'h3CF0;
            14'h116 : data_reg <= 16'h3D2B;
            14'h117 : data_reg <= 16'h092C;
            14'h118 : data_reg <= 16'h213C;
            14'h119 : data_reg <= 16'h2C0B;
            14'h11A : data_reg <= 16'h223C;
            14'h11B : data_reg <= 16'h2C0B;
            14'h11C : data_reg <= 16'h233C;
            14'h11D : data_reg <= 16'h2C0B;
            14'h11E : data_reg <= 16'h243C;
            14'h11F : data_reg <= 16'h2C0B;
            14'h120 : data_reg <= 16'h253C;
            14'h121 : data_reg <= 16'h2C0B;
            14'h122 : data_reg <= 16'h263C;
            14'h123 : data_reg <= 16'h2C0B;
            14'h124 : data_reg <= 16'h273C;
            14'h125 : data_reg <= 16'h2C0B;
            14'h126 : data_reg <= 16'h283C;
            14'h127 : data_reg <= 16'h2C0B;
            14'h128 : data_reg <= 16'h2D3C;
            14'h129 : data_reg <= 16'h2C38;
            14'h12A : data_reg <= 16'h3D16;
            14'h12B : data_reg <= 16'h223C;
            14'h12C : data_reg <= 16'h2C33;
            14'h12D : data_reg <= 16'h2D3C;
            14'h12E : data_reg <= 16'h2C3B;
            14'h12F : data_reg <= 16'h3D10;
            14'h130 : data_reg <= 16'h3C12;
            14'h131 : data_reg <= 16'h4C12;
            14'h132 : data_reg <= 16'h3E4E;
            14'h133 : data_reg <= 16'h02BA;
            14'h134 : data_reg <= 16'h4C13;
            14'h135 : data_reg <= 16'h4E08;
            14'h136 : data_reg <= 16'h3CF0;
            14'h137 : data_reg <= 16'h3D2B;
            14'h138 : data_reg <= 16'h362C;
            14'h139 : data_reg <= 16'h2D3C;
            14'h13A : data_reg <= 16'h2C3B;
            14'h13B : data_reg <= 16'h3D10;
            14'h13C : data_reg <= 16'h3C12;
            14'h13D : data_reg <= 16'h4C12;
            14'h13E : data_reg <= 16'h3E4E;
            14'h13F : data_reg <= 16'h000A;
            14'h140 : data_reg <= 16'h4C13;
            14'h141 : data_reg <= 16'h4E08;
            14'h142 : data_reg <= 16'h3CF0;
            14'h143 : data_reg <= 16'h3D2B;
            14'h144 : data_reg <= 16'h342C;
            14'h145 : data_reg <= 16'h2D3C;
            14'h146 : data_reg <= 16'h2C3B;
            14'h147 : data_reg <= 16'h3D10;
            14'h148 : data_reg <= 16'h3C12;
            14'h149 : data_reg <= 16'h4C12;
            14'h14A : data_reg <= 16'h3E4E;
            14'h14B : data_reg <= 16'h0030;
            14'h14C : data_reg <= 16'h4C13;
            14'h14D : data_reg <= 16'h4E08;
            14'h14E : data_reg <= 16'h3CF0;
            14'h14F : data_reg <= 16'h3D2B;
            14'h150 : data_reg <= 16'h352C;
            14'h151 : data_reg <= 16'h2D3C;
            14'h152 : data_reg <= 16'h2C3B;
            14'h153 : data_reg <= 16'h3D10;
            14'h154 : data_reg <= 16'h3C12;
            14'h155 : data_reg <= 16'h4C12;
            14'h156 : data_reg <= 16'h3E4E;
            14'h157 : data_reg <= 16'h03F0;
            14'h158 : data_reg <= 16'h4C13;
            14'h159 : data_reg <= 16'h4E08;
            14'h15A : data_reg <= 16'h3CF0;
            14'h15B : data_reg <= 16'h3D2B;
            14'h15C : data_reg <= 16'h372C;
            14'h15D : data_reg <= 16'h243C;
            14'h15E : data_reg <= 16'h2C32;
            14'h15F : data_reg <= 16'h0C27;
            14'h160 : data_reg <= 16'h4522;
            14'h161 : data_reg <= 16'h11E3;
            14'h162 : data_reg <= 16'h3343;
            14'h163 : data_reg <= 16'hC110;
            14'h164 : data_reg <= 16'h0126;
            14'h165 : data_reg <= 16'h1009;
            14'h166 : data_reg <= 16'h3CE3;
            14'h167 : data_reg <= 16'h3D28;
            14'h168 : data_reg <= 16'h3C2C;
            14'h169 : data_reg <= 16'h380A;
            14'h16A : data_reg <= 16'h3C2C;
            14'h16B : data_reg <= 16'h370A;
            14'h16C : data_reg <= 16'h3C2C;
            14'h16D : data_reg <= 16'h360A;
            14'h16E : data_reg <= 16'h3C2C;
            14'h16F : data_reg <= 16'h350A;
            14'h170 : data_reg <= 16'h3C2C;
            14'h171 : data_reg <= 16'h340A;
            14'h172 : data_reg <= 16'h3C2C;
            14'h173 : data_reg <= 16'h330A;
            14'h174 : data_reg <= 16'h3C2C;
            14'h175 : data_reg <= 16'h320A;
            14'h176 : data_reg <= 16'h3C2C;
            14'h177 : data_reg <= 16'h3122;
            14'h178 : data_reg <= 16'h3C2C;
            14'h179 : data_reg <= 16'h3B2D;
            14'h17A : data_reg <= 16'h102C;
            14'h17B : data_reg <= 16'h123D;
            14'h17C : data_reg <= 16'h003C;
            14'h17D : data_reg <= 16'h4C12;
            14'h17E : data_reg <= 16'h3E4E;
            14'h17F : data_reg <= 16'h05AD;
            14'h180 : data_reg <= 16'h4C13;
            14'h181 : data_reg <= 16'h4E08;
            14'h182 : data_reg <= 16'h3CF0;
            14'h183 : data_reg <= 16'h3D2B;
            14'h184 : data_reg <= 16'h0C2C;
            14'h185 : data_reg <= 16'h0A3C;
            14'h186 : data_reg <= 16'h2C31;
            14'h187 : data_reg <= 16'h3C0D;
            14'h188 : data_reg <= 16'h3B2D;
            14'h189 : data_reg <= 16'h102C;
            14'h18A : data_reg <= 16'h123D;
            14'h18B : data_reg <= 16'h003C;
            14'h18C : data_reg <= 16'h4C12;
            14'h18D : data_reg <= 16'h3E4E;
            14'h18E : data_reg <= 16'h0030;
            14'h18F : data_reg <= 16'h4C13;
            14'h190 : data_reg <= 16'h4E08;
            14'h191 : data_reg <= 16'h3CF0;
            14'h192 : data_reg <= 16'h3D2B;
            14'h193 : data_reg <= 16'hE22C;
            14'h194 : data_reg <= 16'h4211;
            14'h195 : data_reg <= 16'h10EC;
            14'h196 : data_reg <= 16'h0DEC;
            14'h197 : data_reg <= 16'h223C;
            14'h198 : data_reg <= 16'h2C0B;
            14'h199 : data_reg <= 16'h2D3C;
            14'h19A : data_reg <= 16'h2C3B;
            14'h19B : data_reg <= 16'h3D10;
            14'h19C : data_reg <= 16'h3C12;
            14'h19D : data_reg <= 16'h4C12;
            14'h19E : data_reg <= 16'h3E4E;
            14'h19F : data_reg <= 16'h0064;
            14'h1A0 : data_reg <= 16'h4C13;
            14'h1A1 : data_reg <= 16'h4E08;
            14'h1A2 : data_reg <= 16'h3CF0;
            14'h1A3 : data_reg <= 16'h3D2B;
            14'h1A4 : data_reg <= 16'h4F2C;
            14'h1A5 : data_reg <= 16'h3C32;
            14'h1A6 : data_reg <= 16'h3B2D;
            14'h1A7 : data_reg <= 16'h102C;
            14'h1A8 : data_reg <= 16'h123D;
            14'h1A9 : data_reg <= 16'h003C;
            14'h1AA : data_reg <= 16'h4C12;
            14'h1AB : data_reg <= 16'h3E4E;
            14'h1AC : data_reg <= 16'h0215;
            14'h1AD : data_reg <= 16'h4C13;
            14'h1AE : data_reg <= 16'h4E08;
            14'h1AF : data_reg <= 16'h3CF0;
            14'h1B0 : data_reg <= 16'h3D2B;
            14'h1B1 : data_reg <= 16'h0C2C;
            14'h1B2 : data_reg <= 16'h213C;
            14'h1B3 : data_reg <= 16'h2C0B;
            14'h1B4 : data_reg <= 16'h223C;
            14'h1B5 : data_reg <= 16'h2C31;
            14'h1B6 : data_reg <= 16'h2D3C;
            14'h1B7 : data_reg <= 16'h2C3B;
            14'h1B8 : data_reg <= 16'h3D10;
            14'h1B9 : data_reg <= 16'h3C12;
            14'h1BA : data_reg <= 16'h4C12;
            14'h1BB : data_reg <= 16'h3E4E;
            14'h1BC : data_reg <= 16'h01CF;
            14'h1BD : data_reg <= 16'h4C13;
            14'h1BE : data_reg <= 16'h4E08;
            14'h1BF : data_reg <= 16'h3CF0;
            14'h1C0 : data_reg <= 16'h3D2B;
            14'h1C1 : data_reg <= 16'h0C2C;
            14'h1C2 : data_reg <= 16'h0A3C;
            14'h1C3 : data_reg <= 16'h2C31;
            14'h1C4 : data_reg <= 16'h0A3C;
            14'h1C5 : data_reg <= 16'h2C32;
            14'h1C6 : data_reg <= 16'h3C0D;
            14'h1C7 : data_reg <= 16'h0B23;
            14'h1C8 : data_reg <= 16'h3C2C;
            14'h1C9 : data_reg <= 16'h0B24;
            14'h1CA : data_reg <= 16'h3C2C;
            14'h1CB : data_reg <= 16'h0B25;
            14'h1CC : data_reg <= 16'h3C2C;
            14'h1CD : data_reg <= 16'h0B26;
            14'h1CE : data_reg <= 16'h102C;
            14'h1CF : data_reg <= 16'h3433;
            14'h1D0 : data_reg <= 16'h2D3C;
            14'h1D1 : data_reg <= 16'h2C3B;
            14'h1D2 : data_reg <= 16'h3D10;
            14'h1D3 : data_reg <= 16'h3C12;
            14'h1D4 : data_reg <= 16'h4C12;
            14'h1D5 : data_reg <= 16'h3E4E;
            14'h1D6 : data_reg <= 16'h03DD;
            14'h1D7 : data_reg <= 16'h4C13;
            14'h1D8 : data_reg <= 16'h4E08;
            14'h1D9 : data_reg <= 16'h3CF0;
            14'h1DA : data_reg <= 16'h3D2B;
            14'h1DB : data_reg <= 16'h352C;
            14'h1DC : data_reg <= 16'h2D3C;
            14'h1DD : data_reg <= 16'h2C3B;
            14'h1DE : data_reg <= 16'h3D10;
            14'h1DF : data_reg <= 16'h3C12;
            14'h1E0 : data_reg <= 16'h4C12;
            14'h1E1 : data_reg <= 16'h3E4E;
            14'h1E2 : data_reg <= 16'h03D1;
            14'h1E3 : data_reg <= 16'h4C13;
            14'h1E4 : data_reg <= 16'h4E08;
            14'h1E5 : data_reg <= 16'h3CF0;
            14'h1E6 : data_reg <= 16'h3D2B;
            14'h1E7 : data_reg <= 16'h362C;
            14'h1E8 : data_reg <= 16'h2410;
            14'h1E9 : data_reg <= 16'h25C2;
            14'h1EA : data_reg <= 16'h1109;
            14'h1EB : data_reg <= 16'h3444;
            14'h1EC : data_reg <= 16'h4321;
            14'h1ED : data_reg <= 16'h2633;
            14'h1EE : data_reg <= 16'h233E;
            14'h1EF : data_reg <= 16'h3C31;
            14'h1F0 : data_reg <= 16'h360A;
            14'h1F1 : data_reg <= 16'h3C2C;
            14'h1F2 : data_reg <= 16'h350A;
            14'h1F3 : data_reg <= 16'h3C2C;
            14'h1F4 : data_reg <= 16'h340A;
            14'h1F5 : data_reg <= 16'h3C2C;
            14'h1F6 : data_reg <= 16'h330A;
            14'h1F7 : data_reg <= 16'h0D2C;
            14'h1F8 : data_reg <= 16'h233C;
            14'h1F9 : data_reg <= 16'h2C0B;
            14'h1FA : data_reg <= 16'h253C;
            14'h1FB : data_reg <= 16'h2C0B;
            14'h1FC : data_reg <= 16'h263C;
            14'h1FD : data_reg <= 16'h2C0B;
            14'h1FE : data_reg <= 16'h2D3C;
            14'h1FF : data_reg <= 16'h2C3B;
            14'h200 : data_reg <= 16'h3D10;
            14'h201 : data_reg <= 16'h3C12;
            14'h202 : data_reg <= 16'h4C12;
            14'h203 : data_reg <= 16'h3E4E;
            14'h204 : data_reg <= 16'h042E;
            14'h205 : data_reg <= 16'h4C13;
            14'h206 : data_reg <= 16'h4E08;
            14'h207 : data_reg <= 16'h3CF0;
            14'h208 : data_reg <= 16'h3D2B;
            14'h209 : data_reg <= 16'h352C;
            14'h20A : data_reg <= 16'h2D3C;
            14'h20B : data_reg <= 16'h2C3B;
            14'h20C : data_reg <= 16'h3D10;
            14'h20D : data_reg <= 16'h3C12;
            14'h20E : data_reg <= 16'h4C12;
            14'h20F : data_reg <= 16'h3E4E;
            14'h210 : data_reg <= 16'h043A;
            14'h211 : data_reg <= 16'h4C13;
            14'h212 : data_reg <= 16'h4E08;
            14'h213 : data_reg <= 16'h3CF0;
            14'h214 : data_reg <= 16'h3D2B;
            14'h215 : data_reg <= 16'h362C;
            14'h216 : data_reg <= 16'h3310;
            14'h217 : data_reg <= 16'hD221;
            14'h218 : data_reg <= 16'h0926;
            14'h219 : data_reg <= 16'h5221;
            14'h21A : data_reg <= 16'h1131;
            14'h21B : data_reg <= 16'h3343;
            14'h21C : data_reg <= 16'h3E25;
            14'h21D : data_reg <= 16'h3221;
            14'h21E : data_reg <= 16'h3123;
            14'h21F : data_reg <= 16'h0A3C;
            14'h220 : data_reg <= 16'h2C36;
            14'h221 : data_reg <= 16'h0A3C;
            14'h222 : data_reg <= 16'h2C35;
            14'h223 : data_reg <= 16'h0A3C;
            14'h224 : data_reg <= 16'h2C33;
            14'h225 : data_reg <= 16'h3C0D;
            14'h226 : data_reg <= 16'h0B23;
            14'h227 : data_reg <= 16'h3C2C;
            14'h228 : data_reg <= 16'h0B24;
            14'h229 : data_reg <= 16'h3C2C;
            14'h22A : data_reg <= 16'h0B25;
            14'h22B : data_reg <= 16'h3C2C;
            14'h22C : data_reg <= 16'h0B26;
            14'h22D : data_reg <= 16'h3C2C;
            14'h22E : data_reg <= 16'h0B27;
            14'h22F : data_reg <= 16'h3C2C;
            14'h230 : data_reg <= 16'h3B2D;
            14'h231 : data_reg <= 16'h102C;
            14'h232 : data_reg <= 16'h123D;
            14'h233 : data_reg <= 16'h003C;
            14'h234 : data_reg <= 16'h4C12;
            14'h235 : data_reg <= 16'h3E4E;
            14'h236 : data_reg <= 16'h04CB;
            14'h237 : data_reg <= 16'h4C13;
            14'h238 : data_reg <= 16'h4E08;
            14'h239 : data_reg <= 16'h3CF0;
            14'h23A : data_reg <= 16'h3D2B;
            14'h23B : data_reg <= 16'h352C;
            14'h23C : data_reg <= 16'h2D3C;
            14'h23D : data_reg <= 16'h2C3B;
            14'h23E : data_reg <= 16'h3D10;
            14'h23F : data_reg <= 16'h3C12;
            14'h240 : data_reg <= 16'h4C12;
            14'h241 : data_reg <= 16'h3E4E;
            14'h242 : data_reg <= 16'h04AC;
            14'h243 : data_reg <= 16'h4C13;
            14'h244 : data_reg <= 16'h4E08;
            14'h245 : data_reg <= 16'h3CF0;
            14'h246 : data_reg <= 16'h3D2B;
            14'h247 : data_reg <= 16'h362C;
            14'h248 : data_reg <= 16'h2D3C;
            14'h249 : data_reg <= 16'h2C3B;
            14'h24A : data_reg <= 16'h3D10;
            14'h24B : data_reg <= 16'h3C12;
            14'h24C : data_reg <= 16'h4C12;
            14'h24D : data_reg <= 16'h3E4E;
            14'h24E : data_reg <= 16'h038D;
            14'h24F : data_reg <= 16'h4C13;
            14'h250 : data_reg <= 16'h4E08;
            14'h251 : data_reg <= 16'h3CF0;
            14'h252 : data_reg <= 16'h3D2B;
            14'h253 : data_reg <= 16'h372C;
            14'h254 : data_reg <= 16'h3311;
            14'h255 : data_reg <= 16'h3410;
            14'h256 : data_reg <= 16'hC224;
            14'h257 : data_reg <= 16'h0925;
            14'h258 : data_reg <= 16'h4411;
            14'h259 : data_reg <= 16'h3C34;
            14'h25A : data_reg <= 16'h0B21;
            14'h25B : data_reg <= 16'h3C2C;
            14'h25C : data_reg <= 16'h0B22;
            14'h25D : data_reg <= 16'h232C;
            14'h25E : data_reg <= 16'h2732;
            14'h25F : data_reg <= 16'h210C;
            14'h260 : data_reg <= 16'h3C33;
            14'h261 : data_reg <= 16'h320A;
            14'h262 : data_reg <= 16'h3C2C;
            14'h263 : data_reg <= 16'h310A;
            14'h264 : data_reg <= 16'h262C;
            14'h265 : data_reg <= 16'h233E;
            14'h266 : data_reg <= 16'h3C31;
            14'h267 : data_reg <= 16'h370A;
            14'h268 : data_reg <= 16'h3C2C;
            14'h269 : data_reg <= 16'h360A;
            14'h26A : data_reg <= 16'h3C2C;
            14'h26B : data_reg <= 16'h350A;
            14'h26C : data_reg <= 16'h3C2C;
            14'h26D : data_reg <= 16'h340A;
            14'h26E : data_reg <= 16'h3C2C;
            14'h26F : data_reg <= 16'h330A;
            14'h270 : data_reg <= 16'h0D2C;
            14'h271 : data_reg <= 16'h223C;
            14'h272 : data_reg <= 16'h2C0B;
            14'h273 : data_reg <= 16'h233C;
            14'h274 : data_reg <= 16'h2C0B;
            14'h275 : data_reg <= 16'h243C;
            14'h276 : data_reg <= 16'h2C0B;
            14'h277 : data_reg <= 16'h253C;
            14'h278 : data_reg <= 16'h2C0B;
            14'h279 : data_reg <= 16'h352D;
            14'h27A : data_reg <= 16'h3D16;
            14'h27B : data_reg <= 16'h3221;
            14'h27C : data_reg <= 16'h2D3C;
            14'h27D : data_reg <= 16'h2C3B;
            14'h27E : data_reg <= 16'h3D10;
            14'h27F : data_reg <= 16'h3C12;
            14'h280 : data_reg <= 16'h4C12;
            14'h281 : data_reg <= 16'h3E4E;
            14'h282 : data_reg <= 16'h0512;
            14'h283 : data_reg <= 16'h4C13;
            14'h284 : data_reg <= 16'h4E08;
            14'h285 : data_reg <= 16'h3CF0;
            14'h286 : data_reg <= 16'h3D2B;
            14'h287 : data_reg <= 16'h332C;
            14'h288 : data_reg <= 16'h3410;
            14'h289 : data_reg <= 16'hC4F2;
            14'h28A : data_reg <= 16'h1101;
            14'h28B : data_reg <= 16'h3242;
            14'h28C : data_reg <= 16'h0923;
            14'h28D : data_reg <= 16'h3311;
            14'h28E : data_reg <= 16'h5322;
            14'h28F : data_reg <= 16'h3151;
            14'h290 : data_reg <= 16'h3D25;
            14'h291 : data_reg <= 16'h0A3C;
            14'h292 : data_reg <= 16'h2C35;
            14'h293 : data_reg <= 16'h0A3C;
            14'h294 : data_reg <= 16'h2C34;
            14'h295 : data_reg <= 16'h0A3C;
            14'h296 : data_reg <= 16'h2C33;
            14'h297 : data_reg <= 16'h0A3C;
            14'h298 : data_reg <= 16'h2C32;
            14'h299 : data_reg <= 16'h3C0D;
            14'h29A : data_reg <= 16'h0B21;
            14'h29B : data_reg <= 16'h3C2C;
            14'h29C : data_reg <= 16'h0B22;
            14'h29D : data_reg <= 16'h3C2C;
            14'h29E : data_reg <= 16'h0B23;
            14'h29F : data_reg <= 16'h3C2C;
            14'h2A0 : data_reg <= 16'h0B25;
            14'h2A1 : data_reg <= 16'h3C2C;
            14'h2A2 : data_reg <= 16'h0B26;
            14'h2A3 : data_reg <= 16'h3C2C;
            14'h2A4 : data_reg <= 16'h0B24;
            14'h2A5 : data_reg <= 16'h3C2C;
            14'h2A6 : data_reg <= 16'h342D;
            14'h2A7 : data_reg <= 16'h162C;
            14'h2A8 : data_reg <= 16'h3C3D;
            14'h2A9 : data_reg <= 16'h3B2D;
            14'h2AA : data_reg <= 16'h102C;
            14'h2AB : data_reg <= 16'h123D;
            14'h2AC : data_reg <= 16'h003C;
            14'h2AD : data_reg <= 16'h4C12;
            14'h2AE : data_reg <= 16'h3E4E;
            14'h2AF : data_reg <= 16'h0584;
            14'h2B0 : data_reg <= 16'h4C13;
            14'h2B1 : data_reg <= 16'h4E08;
            14'h2B2 : data_reg <= 16'h3CF0;
            14'h2B3 : data_reg <= 16'h3D2B;
            14'h2B4 : data_reg <= 16'h352C;
            14'h2B5 : data_reg <= 16'h2D3C;
            14'h2B6 : data_reg <= 16'h2C3B;
            14'h2B7 : data_reg <= 16'h3D10;
            14'h2B8 : data_reg <= 16'h3C12;
            14'h2B9 : data_reg <= 16'h4C12;
            14'h2BA : data_reg <= 16'h3E4E;
            14'h2BB : data_reg <= 16'h0592;
            14'h2BC : data_reg <= 16'h4C13;
            14'h2BD : data_reg <= 16'h4E08;
            14'h2BE : data_reg <= 16'h3CF0;
            14'h2BF : data_reg <= 16'h3D2B;
            14'h2C0 : data_reg <= 16'h362C;
            14'h2C1 : data_reg <= 16'h3C11;
            14'h2C2 : data_reg <= 16'hC210;
            14'h2C3 : data_reg <= 16'h0926;
            14'h2C4 : data_reg <= 16'hE123;
            14'h2C5 : data_reg <= 16'h4C21;
            14'h2C6 : data_reg <= 16'h2231;
            14'h2C7 : data_reg <= 16'h325C;
            14'h2C8 : data_reg <= 16'h3E25;
            14'h2C9 : data_reg <= 16'h3D24;
            14'h2CA : data_reg <= 16'h0A3C;
            14'h2CB : data_reg <= 16'h2C34;
            14'h2CC : data_reg <= 16'h0A3C;
            14'h2CD : data_reg <= 16'h2C36;
            14'h2CE : data_reg <= 16'h0A3C;
            14'h2CF : data_reg <= 16'h2C34;
            14'h2D0 : data_reg <= 16'h0A3C;
            14'h2D1 : data_reg <= 16'h2C33;
            14'h2D2 : data_reg <= 16'h0A3C;
            14'h2D3 : data_reg <= 16'h2C32;
            14'h2D4 : data_reg <= 16'h0A3C;
            14'h2D5 : data_reg <= 16'h2C31;
            14'h2D6 : data_reg <= 16'h3C0D;
            14'h2D7 : data_reg <= 16'h0B22;
            14'h2D8 : data_reg <= 16'h3C2C;
            14'h2D9 : data_reg <= 16'h0B23;
            14'h2DA : data_reg <= 16'h3C2C;
            14'h2DB : data_reg <= 16'h0B24;
            14'h2DC : data_reg <= 16'h3C2C;
            14'h2DD : data_reg <= 16'h0B25;
            14'h2DE : data_reg <= 16'h3C2C;
            14'h2DF : data_reg <= 16'h0B26;
            14'h2E0 : data_reg <= 16'h3C2C;
            14'h2E1 : data_reg <= 16'h0B27;
            14'h2E2 : data_reg <= 16'h3C2C;
            14'h2E3 : data_reg <= 16'h0B28;
            14'h2E4 : data_reg <= 16'h3C2C;
            14'h2E5 : data_reg <= 16'h0B21;
            14'h2E6 : data_reg <= 16'h3C2C;
            14'h2E7 : data_reg <= 16'h3B2D;
            14'h2E8 : data_reg <= 16'h102C;
            14'h2E9 : data_reg <= 16'h123D;
            14'h2EA : data_reg <= 16'h003C;
            14'h2EB : data_reg <= 16'h4C12;
            14'h2EC : data_reg <= 16'h3E4E;
            14'h2ED : data_reg <= 16'h04E2;
            14'h2EE : data_reg <= 16'h4C13;
            14'h2EF : data_reg <= 16'h4E08;
            14'h2F0 : data_reg <= 16'h3CF0;
            14'h2F1 : data_reg <= 16'h3D2B;
            14'h2F2 : data_reg <= 16'h0C2C;
            14'h2F3 : data_reg <= 16'h3221;
            14'h2F4 : data_reg <= 16'h0A3C;
            14'h2F5 : data_reg <= 16'h2C31;
            14'h2F6 : data_reg <= 16'h3310;
            14'h2F7 : data_reg <= 16'h3C11;
            14'h2F8 : data_reg <= 16'hBC22;
            14'h2F9 : data_reg <= 16'h3C34;
            14'h2FA : data_reg <= 16'h3B2D;
            14'h2FB : data_reg <= 16'h102C;
            14'h2FC : data_reg <= 16'h123D;
            14'h2FD : data_reg <= 16'h003C;
            14'h2FE : data_reg <= 16'h4C12;
            14'h2FF : data_reg <= 16'h3E4E;
            14'h300 : data_reg <= 16'h062A;
            14'h301 : data_reg <= 16'h4C13;
            14'h302 : data_reg <= 16'h4E08;
            14'h303 : data_reg <= 16'h3CF0;
            14'h304 : data_reg <= 16'h3D2B;
            14'h305 : data_reg <= 16'h352C;
            14'h306 : data_reg <= 16'h2D3C;
            14'h307 : data_reg <= 16'h2C3B;
            14'h308 : data_reg <= 16'h3D10;
            14'h309 : data_reg <= 16'h3C12;
            14'h30A : data_reg <= 16'h4C12;
            14'h30B : data_reg <= 16'h3E4E;
            14'h30C : data_reg <= 16'h0645;
            14'h30D : data_reg <= 16'h4C13;
            14'h30E : data_reg <= 16'h4E08;
            14'h30F : data_reg <= 16'h3CF0;
            14'h310 : data_reg <= 16'h3D2B;
            14'h311 : data_reg <= 16'h362C;
            14'h312 : data_reg <= 16'h2D3C;
            14'h313 : data_reg <= 16'h2C37;
            14'h314 : data_reg <= 16'h3D16;
            14'h315 : data_reg <= 16'hC423;
            14'h316 : data_reg <= 16'h0926;
            14'h317 : data_reg <= 16'h4321;
            14'h318 : data_reg <= 16'hF03B;
            14'h319 : data_reg <= 16'h110B;
            14'h31A : data_reg <= 16'h213C;
            14'h31B : data_reg <= 16'h5342;
            14'h31C : data_reg <= 16'h3C5C;
            14'h31D : data_reg <= 16'h38FC;
            14'h31E : data_reg <= 16'hEC0A;
            14'h31F : data_reg <= 16'hEB28;
            14'h320 : data_reg <= 16'h4311;
            14'h321 : data_reg <= 16'h2533;
            14'h322 : data_reg <= 16'h273E;
            14'h323 : data_reg <= 16'h3C3D;
            14'h324 : data_reg <= 16'h380A;
            14'h325 : data_reg <= 16'h3C2C;
            14'h326 : data_reg <= 16'h370A;
            14'h327 : data_reg <= 16'h3C2C;
            14'h328 : data_reg <= 16'h360A;
            14'h329 : data_reg <= 16'h3C2C;
            14'h32A : data_reg <= 16'h350A;
            14'h32B : data_reg <= 16'h3C2C;
            14'h32C : data_reg <= 16'h340A;
            14'h32D : data_reg <= 16'h3C2C;
            14'h32E : data_reg <= 16'h330A;
            14'h32F : data_reg <= 16'h3C2C;
            14'h330 : data_reg <= 16'h320A;
            14'h331 : data_reg <= 16'h0D2C;
            14'h332 : data_reg <= 16'h6548;
            14'h333 : data_reg <= 16'h6C6C;
            14'h334 : data_reg <= 16'h2C6F;
            14'h335 : data_reg <= 16'h7720;
            14'h336 : data_reg <= 16'h726F;
            14'h337 : data_reg <= 16'h646C;
            14'h338 : data_reg <= 16'h0D21;
            14'h339 : data_reg <= 16'h000A;
            14'h33A : data_reg <= 16'h2D3C;
            14'h33B : data_reg <= 16'h2C3B;
            14'h33C : data_reg <= 16'h3D10;
            14'h33D : data_reg <= 16'h3C12;
            14'h33E : data_reg <= 16'h4C12;
            14'h33F : data_reg <= 16'h3E4E;
            14'h340 : data_reg <= 16'h0664;
            14'h341 : data_reg <= 16'h4C13;
            14'h342 : data_reg <= 16'h4E08;
            14'h343 : data_reg <= 16'h3CF0;
            14'h344 : data_reg <= 16'h3D2B;
            14'h345 : data_reg <= 16'h312C;
            14'h346 : data_reg <= 16'h2D3C;
            14'h347 : data_reg <= 16'h2C3B;
            14'h348 : data_reg <= 16'h3D10;
            14'h349 : data_reg <= 16'h3C12;
            14'h34A : data_reg <= 16'h4C12;
            14'h34B : data_reg <= 16'h3E4E;
            14'h34C : data_reg <= 16'h01CF;
            14'h34D : data_reg <= 16'h4C13;
            14'h34E : data_reg <= 16'h4E08;
            14'h34F : data_reg <= 16'h3CF0;
            14'h350 : data_reg <= 16'h3D2B;
            14'h351 : data_reg <= 16'h0C2C;
            14'h352 : data_reg <= 16'h000E;
            default : data_reg <= 0;
        endcase
    assign data = ( enable ? data_reg : 0 );
endmodule
