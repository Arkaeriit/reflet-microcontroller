//The code used to make this ROM is in software/helloWorld.asm
module rom2(input clk, input enable, input [10-1:0] addr, output [16-1:0] data_out);
    reg [16-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            10'h0 : data_reg <= 16'h5341;
            10'h1 : data_reg <= 16'h4D52;
            10'h2 : data_reg <= 16'h3C3C;
            10'h3 : data_reg <= 16'h3B2D;
            10'h4 : data_reg <= 16'h102C;
            10'h5 : data_reg <= 16'h003D;
            10'h6 : data_reg <= 16'h0000;
            10'h7 : data_reg <= 16'h3C12;
            10'h8 : data_reg <= 16'h4C12;
            10'h9 : data_reg <= 16'h3E4E;
            10'hA : data_reg <= 16'h8000;
            10'hB : data_reg <= 16'h4C13;
            10'hC : data_reg <= 16'h4E08;
            10'hD : data_reg <= 16'h3CF0;
            10'hE : data_reg <= 16'h3D2B;
            10'hF : data_reg <= 16'h3F2C;
            10'h10 : data_reg <= 16'h3C2C;
            10'h11 : data_reg <= 16'h3B2D;
            10'h12 : data_reg <= 16'h102C;
            10'h13 : data_reg <= 16'h003D;
            10'h14 : data_reg <= 16'h0000;
            10'h15 : data_reg <= 16'h3C12;
            10'h16 : data_reg <= 16'h4C12;
            10'h17 : data_reg <= 16'h3E4E;
            10'h18 : data_reg <= 16'h0668;
            10'h19 : data_reg <= 16'h4C13;
            10'h1A : data_reg <= 16'h4E08;
            10'h1B : data_reg <= 16'h3CF0;
            10'h1C : data_reg <= 16'h3D2B;
            10'h1D : data_reg <= 16'h3E2C;
            10'h1E : data_reg <= 16'h223C;
            10'h1F : data_reg <= 16'h2C0B;
            10'h20 : data_reg <= 16'h243C;
            10'h21 : data_reg <= 16'h2C0B;
            10'h22 : data_reg <= 16'h2D3C;
            10'h23 : data_reg <= 16'h2C3B;
            10'h24 : data_reg <= 16'h3D10;
            10'h25 : data_reg <= 16'h0000;
            10'h26 : data_reg <= 16'h3C12;
            10'h27 : data_reg <= 16'h4C12;
            10'h28 : data_reg <= 16'h3E4E;
            10'h29 : data_reg <= 16'h00E0;
            10'h2A : data_reg <= 16'h4C13;
            10'h2B : data_reg <= 16'h4E08;
            10'h2C : data_reg <= 16'h3CF0;
            10'h2D : data_reg <= 16'h3D2B;
            10'h2E : data_reg <= 16'hF02C;
            10'h2F : data_reg <= 16'h3203;
            10'h30 : data_reg <= 16'h2D3C;
            10'h31 : data_reg <= 16'h2C3B;
            10'h32 : data_reg <= 16'h3D10;
            10'h33 : data_reg <= 16'h0000;
            10'h34 : data_reg <= 16'h3C12;
            10'h35 : data_reg <= 16'h4C12;
            10'h36 : data_reg <= 16'h3E4E;
            10'h37 : data_reg <= 16'h007A;
            10'h38 : data_reg <= 16'h4C13;
            10'h39 : data_reg <= 16'h4E08;
            10'h3A : data_reg <= 16'h3CF0;
            10'h3B : data_reg <= 16'h3D2B;
            10'h3C : data_reg <= 16'h342C;
            10'h3D : data_reg <= 16'h3CF2;
            10'h3E : data_reg <= 16'hCC10;
            10'h3F : data_reg <= 16'h0924;
            10'h40 : data_reg <= 16'h4211;
            10'h41 : data_reg <= 16'h213C;
            10'h42 : data_reg <= 16'h10EC;
            10'h43 : data_reg <= 16'h03E2;
            10'h44 : data_reg <= 16'h0A3C;
            10'h45 : data_reg <= 16'h2C34;
            10'h46 : data_reg <= 16'h0A3C;
            10'h47 : data_reg <= 16'h2C32;
            10'h48 : data_reg <= 16'h3C0D;
            10'h49 : data_reg <= 16'h0B21;
            10'h4A : data_reg <= 16'h1A2C;
            10'h4B : data_reg <= 16'h3C31;
            10'h4C : data_reg <= 16'h3B2D;
            10'h4D : data_reg <= 16'h102C;
            10'h4E : data_reg <= 16'h003D;
            10'h4F : data_reg <= 16'h0000;
            10'h50 : data_reg <= 16'h3C12;
            10'h51 : data_reg <= 16'h4C12;
            10'h52 : data_reg <= 16'h3E4E;
            10'h53 : data_reg <= 16'h003C;
            10'h54 : data_reg <= 16'h4C13;
            10'h55 : data_reg <= 16'h4E08;
            10'h56 : data_reg <= 16'h3CF0;
            10'h57 : data_reg <= 16'h3D2B;
            10'h58 : data_reg <= 16'h0C2C;
            10'h59 : data_reg <= 16'h311D;
            10'h5A : data_reg <= 16'h2D3C;
            10'h5B : data_reg <= 16'h2C3B;
            10'h5C : data_reg <= 16'h3D10;
            10'h5D : data_reg <= 16'h0000;
            10'h5E : data_reg <= 16'h3C12;
            10'h5F : data_reg <= 16'h4C12;
            10'h60 : data_reg <= 16'h3E4E;
            10'h61 : data_reg <= 16'h003C;
            10'h62 : data_reg <= 16'h4C13;
            10'h63 : data_reg <= 16'h4E08;
            10'h64 : data_reg <= 16'h3CF0;
            10'h65 : data_reg <= 16'h3D2B;
            10'h66 : data_reg <= 16'h0C2C;
            10'h67 : data_reg <= 16'h0A3C;
            10'h68 : data_reg <= 16'h2C31;
            10'h69 : data_reg <= 16'h000D;
            10'h6A : data_reg <= 16'h8000;
            10'h6B : data_reg <= 16'hFF00;
            10'h6C : data_reg <= 16'hFF04;
            10'h6D : data_reg <= 16'hFF08;
            10'h6E : data_reg <= 16'hFF10;
            10'h6F : data_reg <= 16'hFF13;
            10'h70 : data_reg <= 16'hFF16;
            10'h71 : data_reg <= 16'hFF1A;
            10'h72 : data_reg <= 16'hFF1C;
            10'h73 : data_reg <= 16'hFF1F;
            10'h74 : data_reg <= 16'hFF21;
            10'h75 : data_reg <= 16'hFF22;
            10'h76 : data_reg <= 16'h213C;
            10'h77 : data_reg <= 16'h2C0B;
            10'h78 : data_reg <= 16'h223C;
            10'h79 : data_reg <= 16'h2C0B;
            10'h7A : data_reg <= 16'h233C;
            10'h7B : data_reg <= 16'h2C0B;
            10'h7C : data_reg <= 16'h243C;
            10'h7D : data_reg <= 16'h2C0B;
            10'h7E : data_reg <= 16'h253C;
            10'h7F : data_reg <= 16'h2C0B;
            10'h80 : data_reg <= 16'h263C;
            10'h81 : data_reg <= 16'h2C0B;
            10'h82 : data_reg <= 16'h2D3C;
            10'h83 : data_reg <= 16'h2C3B;
            10'h84 : data_reg <= 16'h3D10;
            10'h85 : data_reg <= 16'h0000;
            10'h86 : data_reg <= 16'h3C12;
            10'h87 : data_reg <= 16'h4C12;
            10'h88 : data_reg <= 16'h3E4E;
            10'h89 : data_reg <= 16'h0154;
            10'h8A : data_reg <= 16'h4C13;
            10'h8B : data_reg <= 16'h4E08;
            10'h8C : data_reg <= 16'h3CF0;
            10'h8D : data_reg <= 16'h3D2B;
            10'h8E : data_reg <= 16'h332C;
            10'h8F : data_reg <= 16'h2D3C;
            10'h90 : data_reg <= 16'h2C3B;
            10'h91 : data_reg <= 16'h3D10;
            10'h92 : data_reg <= 16'h0000;
            10'h93 : data_reg <= 16'h3C12;
            10'h94 : data_reg <= 16'h4C12;
            10'h95 : data_reg <= 16'h3E4E;
            10'h96 : data_reg <= 16'h0172;
            10'h97 : data_reg <= 16'h4C13;
            10'h98 : data_reg <= 16'h4E08;
            10'h99 : data_reg <= 16'h3CF0;
            10'h9A : data_reg <= 16'h3D2B;
            10'h9B : data_reg <= 16'h342C;
            10'h9C : data_reg <= 16'h3511;
            10'h9D : data_reg <= 16'h2D3C;
            10'h9E : data_reg <= 16'h2C3B;
            10'h9F : data_reg <= 16'h3D10;
            10'hA0 : data_reg <= 16'h0000;
            10'hA1 : data_reg <= 16'h3C12;
            10'hA2 : data_reg <= 16'h4C12;
            10'hA3 : data_reg <= 16'h3E4E;
            10'hA4 : data_reg <= 16'h003C;
            10'hA5 : data_reg <= 16'h4C13;
            10'hA6 : data_reg <= 16'h4E08;
            10'hA7 : data_reg <= 16'h3CF0;
            10'hA8 : data_reg <= 16'h3D2B;
            10'hA9 : data_reg <= 16'h362C;
            10'hAA : data_reg <= 16'hC210;
            10'hAB : data_reg <= 16'h0924;
            10'hAC : data_reg <= 16'hF103;
            10'hAD : data_reg <= 16'h3C03;
            10'hAE : data_reg <= 16'h213C;
            10'hAF : data_reg <= 16'h2C0B;
            10'hB0 : data_reg <= 16'h2C3C;
            10'hB1 : data_reg <= 16'h2C31;
            10'hB2 : data_reg <= 16'h0C26;
            10'hB3 : data_reg <= 16'h0A3C;
            10'hB4 : data_reg <= 16'h2C31;
            10'hB5 : data_reg <= 16'h4521;
            10'hB6 : data_reg <= 16'h2231;
            10'hB7 : data_reg <= 16'h3255;
            10'hB8 : data_reg <= 16'h3E23;
            10'hB9 : data_reg <= 16'h0A3C;
            10'hBA : data_reg <= 16'h2C36;
            10'hBB : data_reg <= 16'h0A3C;
            10'hBC : data_reg <= 16'h2C35;
            10'hBD : data_reg <= 16'h0A3C;
            10'hBE : data_reg <= 16'h2C34;
            10'hBF : data_reg <= 16'h0A3C;
            10'hC0 : data_reg <= 16'h2C33;
            10'hC1 : data_reg <= 16'h0A3C;
            10'hC2 : data_reg <= 16'h2C32;
            10'hC3 : data_reg <= 16'h0A3C;
            10'hC4 : data_reg <= 16'h2C31;
            10'hC5 : data_reg <= 16'h3C0D;
            10'hC6 : data_reg <= 16'h0B22;
            10'hC7 : data_reg <= 16'h3C2C;
            10'hC8 : data_reg <= 16'h0B21;
            10'hC9 : data_reg <= 16'h3C2C;
            10'hCA : data_reg <= 16'h3B2D;
            10'hCB : data_reg <= 16'h102C;
            10'hCC : data_reg <= 16'h003D;
            10'hCD : data_reg <= 16'h0000;
            10'hCE : data_reg <= 16'h3C12;
            10'hCF : data_reg <= 16'h4C12;
            10'hD0 : data_reg <= 16'h3E4E;
            10'hD1 : data_reg <= 16'h04CA;
            10'hD2 : data_reg <= 16'h4C13;
            10'hD3 : data_reg <= 16'h4E08;
            10'hD4 : data_reg <= 16'h3CF0;
            10'hD5 : data_reg <= 16'h3D2B;
            10'hD6 : data_reg <= 16'h0C2C;
            10'hD7 : data_reg <= 16'h213C;
            10'hD8 : data_reg <= 16'h2C32;
            10'hD9 : data_reg <= 16'h0A3C;
            10'hDA : data_reg <= 16'h2C31;
            10'hDB : data_reg <= 16'h2D3C;
            10'hDC : data_reg <= 16'h2C3B;
            10'hDD : data_reg <= 16'h3D10;
            10'hDE : data_reg <= 16'h0000;
            10'hDF : data_reg <= 16'h3C12;
            10'hE0 : data_reg <= 16'h4C12;
            10'hE1 : data_reg <= 16'h3E4E;
            10'hE2 : data_reg <= 16'h00EC;
            10'hE3 : data_reg <= 16'h4C13;
            10'hE4 : data_reg <= 16'h4E08;
            10'hE5 : data_reg <= 16'h3CF0;
            10'hE6 : data_reg <= 16'h3D2B;
            10'hE7 : data_reg <= 16'h0C2C;
            10'hE8 : data_reg <= 16'h0A3C;
            10'hE9 : data_reg <= 16'h2C32;
            10'hEA : data_reg <= 16'h100D;
            10'hEB : data_reg <= 16'h3CC1;
            10'hEC : data_reg <= 16'h3B2D;
            10'hED : data_reg <= 16'h102C;
            10'hEE : data_reg <= 16'h003D;
            10'hEF : data_reg <= 16'h0000;
            10'hF0 : data_reg <= 16'h3C12;
            10'hF1 : data_reg <= 16'h4C12;
            10'hF2 : data_reg <= 16'h3E4E;
            10'hF3 : data_reg <= 16'h02E1;
            10'hF4 : data_reg <= 16'h4C13;
            10'hF5 : data_reg <= 16'h4E08;
            10'hF6 : data_reg <= 16'h3CF0;
            10'hF7 : data_reg <= 16'h3D2B;
            10'hF8 : data_reg <= 16'h092C;
            10'hF9 : data_reg <= 16'h213C;
            10'hFA : data_reg <= 16'h2C0B;
            10'hFB : data_reg <= 16'h223C;
            10'hFC : data_reg <= 16'h2C0B;
            10'hFD : data_reg <= 16'h233C;
            10'hFE : data_reg <= 16'h2C0B;
            10'hFF : data_reg <= 16'h243C;
            10'h100 : data_reg <= 16'h2C0B;
            10'h101 : data_reg <= 16'h253C;
            10'h102 : data_reg <= 16'h2C0B;
            10'h103 : data_reg <= 16'h263C;
            10'h104 : data_reg <= 16'h2C0B;
            10'h105 : data_reg <= 16'h273C;
            10'h106 : data_reg <= 16'h2C0B;
            10'h107 : data_reg <= 16'h283C;
            10'h108 : data_reg <= 16'h2C0B;
            10'h109 : data_reg <= 16'h2D3C;
            10'h10A : data_reg <= 16'h2C38;
            10'h10B : data_reg <= 16'h3D16;
            10'h10C : data_reg <= 16'h223C;
            10'h10D : data_reg <= 16'h2C33;
            10'h10E : data_reg <= 16'h2D3C;
            10'h10F : data_reg <= 16'h2C3B;
            10'h110 : data_reg <= 16'h3D10;
            10'h111 : data_reg <= 16'h0000;
            10'h112 : data_reg <= 16'h3C12;
            10'h113 : data_reg <= 16'h4C12;
            10'h114 : data_reg <= 16'h3E4E;
            10'h115 : data_reg <= 16'h028A;
            10'h116 : data_reg <= 16'h4C13;
            10'h117 : data_reg <= 16'h4E08;
            10'h118 : data_reg <= 16'h3CF0;
            10'h119 : data_reg <= 16'h3D2B;
            10'h11A : data_reg <= 16'h362C;
            10'h11B : data_reg <= 16'h3C3C;
            10'h11C : data_reg <= 16'h3B2D;
            10'h11D : data_reg <= 16'h102C;
            10'h11E : data_reg <= 16'h003D;
            10'h11F : data_reg <= 16'h0000;
            10'h120 : data_reg <= 16'h3C12;
            10'h121 : data_reg <= 16'h4C12;
            10'h122 : data_reg <= 16'h3E4E;
            10'h123 : data_reg <= 16'h000A;
            10'h124 : data_reg <= 16'h4C13;
            10'h125 : data_reg <= 16'h4E08;
            10'h126 : data_reg <= 16'h3CF0;
            10'h127 : data_reg <= 16'h3D2B;
            10'h128 : data_reg <= 16'h342C;
            10'h129 : data_reg <= 16'h3C2C;
            10'h12A : data_reg <= 16'h2D3C;
            10'h12B : data_reg <= 16'h2C3B;
            10'h12C : data_reg <= 16'h3D10;
            10'h12D : data_reg <= 16'h0000;
            10'h12E : data_reg <= 16'h3C12;
            10'h12F : data_reg <= 16'h4C12;
            10'h130 : data_reg <= 16'h3E4E;
            10'h131 : data_reg <= 16'h0030;
            10'h132 : data_reg <= 16'h4C13;
            10'h133 : data_reg <= 16'h4E08;
            10'h134 : data_reg <= 16'h3CF0;
            10'h135 : data_reg <= 16'h3D2B;
            10'h136 : data_reg <= 16'h352C;
            10'h137 : data_reg <= 16'h3C2C;
            10'h138 : data_reg <= 16'h3B2D;
            10'h139 : data_reg <= 16'h102C;
            10'h13A : data_reg <= 16'h003D;
            10'h13B : data_reg <= 16'h0000;
            10'h13C : data_reg <= 16'h3C12;
            10'h13D : data_reg <= 16'h4C12;
            10'h13E : data_reg <= 16'h3E4E;
            10'h13F : data_reg <= 16'h03CE;
            10'h140 : data_reg <= 16'h4C13;
            10'h141 : data_reg <= 16'h4E08;
            10'h142 : data_reg <= 16'h3CF0;
            10'h143 : data_reg <= 16'h3D2B;
            10'h144 : data_reg <= 16'h372C;
            10'h145 : data_reg <= 16'h243C;
            10'h146 : data_reg <= 16'h2C32;
            10'h147 : data_reg <= 16'h0C27;
            10'h148 : data_reg <= 16'h4522;
            10'h149 : data_reg <= 16'h11E3;
            10'h14A : data_reg <= 16'h3343;
            10'h14B : data_reg <= 16'hC110;
            10'h14C : data_reg <= 16'h0126;
            10'h14D : data_reg <= 16'h1009;
            10'h14E : data_reg <= 16'h3CE3;
            10'h14F : data_reg <= 16'h3D28;
            10'h150 : data_reg <= 16'h3C2C;
            10'h151 : data_reg <= 16'h380A;
            10'h152 : data_reg <= 16'h3C2C;
            10'h153 : data_reg <= 16'h370A;
            10'h154 : data_reg <= 16'h3C2C;
            10'h155 : data_reg <= 16'h360A;
            10'h156 : data_reg <= 16'h3C2C;
            10'h157 : data_reg <= 16'h350A;
            10'h158 : data_reg <= 16'h3C2C;
            10'h159 : data_reg <= 16'h340A;
            10'h15A : data_reg <= 16'h3C2C;
            10'h15B : data_reg <= 16'h330A;
            10'h15C : data_reg <= 16'h3C2C;
            10'h15D : data_reg <= 16'h320A;
            10'h15E : data_reg <= 16'h3C2C;
            10'h15F : data_reg <= 16'h3122;
            10'h160 : data_reg <= 16'h3C2C;
            10'h161 : data_reg <= 16'h3B2D;
            10'h162 : data_reg <= 16'h102C;
            10'h163 : data_reg <= 16'h003D;
            10'h164 : data_reg <= 16'h0000;
            10'h165 : data_reg <= 16'h3C12;
            10'h166 : data_reg <= 16'h4C12;
            10'h167 : data_reg <= 16'h3E4E;
            10'h168 : data_reg <= 16'h059B;
            10'h169 : data_reg <= 16'h4C13;
            10'h16A : data_reg <= 16'h4E08;
            10'h16B : data_reg <= 16'h3CF0;
            10'h16C : data_reg <= 16'h3D2B;
            10'h16D : data_reg <= 16'h0C2C;
            10'h16E : data_reg <= 16'h0A3C;
            10'h16F : data_reg <= 16'h2C31;
            10'h170 : data_reg <= 16'h3C0D;
            10'h171 : data_reg <= 16'h3B2D;
            10'h172 : data_reg <= 16'h102C;
            10'h173 : data_reg <= 16'h003D;
            10'h174 : data_reg <= 16'h0000;
            10'h175 : data_reg <= 16'h3C12;
            10'h176 : data_reg <= 16'h4C12;
            10'h177 : data_reg <= 16'h3E4E;
            10'h178 : data_reg <= 16'h0030;
            10'h179 : data_reg <= 16'h4C13;
            10'h17A : data_reg <= 16'h4E08;
            10'h17B : data_reg <= 16'h3CF0;
            10'h17C : data_reg <= 16'h3D2B;
            10'h17D : data_reg <= 16'hE22C;
            10'h17E : data_reg <= 16'h4211;
            10'h17F : data_reg <= 16'h10EC;
            10'h180 : data_reg <= 16'h0DEC;
            10'h181 : data_reg <= 16'h223C;
            10'h182 : data_reg <= 16'h2C0B;
            10'h183 : data_reg <= 16'h2D3C;
            10'h184 : data_reg <= 16'h2C3B;
            10'h185 : data_reg <= 16'h3D10;
            10'h186 : data_reg <= 16'h0000;
            10'h187 : data_reg <= 16'h3C12;
            10'h188 : data_reg <= 16'h4C12;
            10'h189 : data_reg <= 16'h3E4E;
            10'h18A : data_reg <= 16'h0064;
            10'h18B : data_reg <= 16'h4C13;
            10'h18C : data_reg <= 16'h4E08;
            10'h18D : data_reg <= 16'h3CF0;
            10'h18E : data_reg <= 16'h3D2B;
            10'h18F : data_reg <= 16'h4F2C;
            10'h190 : data_reg <= 16'h3C32;
            10'h191 : data_reg <= 16'h3B2D;
            10'h192 : data_reg <= 16'h102C;
            10'h193 : data_reg <= 16'h003D;
            10'h194 : data_reg <= 16'h0000;
            10'h195 : data_reg <= 16'h3C12;
            10'h196 : data_reg <= 16'h4C12;
            10'h197 : data_reg <= 16'h3E4E;
            10'h198 : data_reg <= 16'h01D5;
            10'h199 : data_reg <= 16'h4C13;
            10'h19A : data_reg <= 16'h4E08;
            10'h19B : data_reg <= 16'h3CF0;
            10'h19C : data_reg <= 16'h3D2B;
            10'h19D : data_reg <= 16'h0C2C;
            10'h19E : data_reg <= 16'h213C;
            10'h19F : data_reg <= 16'h2C0B;
            10'h1A0 : data_reg <= 16'h223C;
            10'h1A1 : data_reg <= 16'h2C31;
            10'h1A2 : data_reg <= 16'h2D3C;
            10'h1A3 : data_reg <= 16'h2C3B;
            10'h1A4 : data_reg <= 16'h3D10;
            10'h1A5 : data_reg <= 16'h0000;
            10'h1A6 : data_reg <= 16'h3C12;
            10'h1A7 : data_reg <= 16'h4C12;
            10'h1A8 : data_reg <= 16'h3E4E;
            10'h1A9 : data_reg <= 16'h018B;
            10'h1AA : data_reg <= 16'h4C13;
            10'h1AB : data_reg <= 16'h4E08;
            10'h1AC : data_reg <= 16'h3CF0;
            10'h1AD : data_reg <= 16'h3D2B;
            10'h1AE : data_reg <= 16'h0C2C;
            10'h1AF : data_reg <= 16'h0A3C;
            10'h1B0 : data_reg <= 16'h2C31;
            10'h1B1 : data_reg <= 16'h0A3C;
            10'h1B2 : data_reg <= 16'h2C32;
            10'h1B3 : data_reg <= 16'h3C0D;
            10'h1B4 : data_reg <= 16'h0B23;
            10'h1B5 : data_reg <= 16'h3C2C;
            10'h1B6 : data_reg <= 16'h0B24;
            10'h1B7 : data_reg <= 16'h3C2C;
            10'h1B8 : data_reg <= 16'h0B25;
            10'h1B9 : data_reg <= 16'h3C2C;
            10'h1BA : data_reg <= 16'h0B26;
            10'h1BB : data_reg <= 16'h102C;
            10'h1BC : data_reg <= 16'h3433;
            10'h1BD : data_reg <= 16'h2D3C;
            10'h1BE : data_reg <= 16'h2C3B;
            10'h1BF : data_reg <= 16'h3D10;
            10'h1C0 : data_reg <= 16'h0000;
            10'h1C1 : data_reg <= 16'h3C12;
            10'h1C2 : data_reg <= 16'h4C12;
            10'h1C3 : data_reg <= 16'h3E4E;
            10'h1C4 : data_reg <= 16'h03BB;
            10'h1C5 : data_reg <= 16'h4C13;
            10'h1C6 : data_reg <= 16'h4E08;
            10'h1C7 : data_reg <= 16'h3CF0;
            10'h1C8 : data_reg <= 16'h3D2B;
            10'h1C9 : data_reg <= 16'h352C;
            10'h1CA : data_reg <= 16'h2D3C;
            10'h1CB : data_reg <= 16'h2C3B;
            10'h1CC : data_reg <= 16'h3D10;
            10'h1CD : data_reg <= 16'h0000;
            10'h1CE : data_reg <= 16'h3C12;
            10'h1CF : data_reg <= 16'h4C12;
            10'h1D0 : data_reg <= 16'h3E4E;
            10'h1D1 : data_reg <= 16'h03AF;
            10'h1D2 : data_reg <= 16'h4C13;
            10'h1D3 : data_reg <= 16'h4E08;
            10'h1D4 : data_reg <= 16'h3CF0;
            10'h1D5 : data_reg <= 16'h3D2B;
            10'h1D6 : data_reg <= 16'h362C;
            10'h1D7 : data_reg <= 16'h2410;
            10'h1D8 : data_reg <= 16'h25C2;
            10'h1D9 : data_reg <= 16'h1109;
            10'h1DA : data_reg <= 16'h3444;
            10'h1DB : data_reg <= 16'h4321;
            10'h1DC : data_reg <= 16'h2633;
            10'h1DD : data_reg <= 16'h233E;
            10'h1DE : data_reg <= 16'h3C31;
            10'h1DF : data_reg <= 16'h360A;
            10'h1E0 : data_reg <= 16'h3C2C;
            10'h1E1 : data_reg <= 16'h350A;
            10'h1E2 : data_reg <= 16'h3C2C;
            10'h1E3 : data_reg <= 16'h340A;
            10'h1E4 : data_reg <= 16'h3C2C;
            10'h1E5 : data_reg <= 16'h330A;
            10'h1E6 : data_reg <= 16'h0D2C;
            10'h1E7 : data_reg <= 16'h233C;
            10'h1E8 : data_reg <= 16'h2C0B;
            10'h1E9 : data_reg <= 16'h253C;
            10'h1EA : data_reg <= 16'h2C0B;
            10'h1EB : data_reg <= 16'h263C;
            10'h1EC : data_reg <= 16'h2C0B;
            10'h1ED : data_reg <= 16'h2D3C;
            10'h1EE : data_reg <= 16'h2C3B;
            10'h1EF : data_reg <= 16'h3D10;
            10'h1F0 : data_reg <= 16'h0000;
            10'h1F1 : data_reg <= 16'h3C12;
            10'h1F2 : data_reg <= 16'h4C12;
            10'h1F3 : data_reg <= 16'h3E4E;
            10'h1F4 : data_reg <= 16'h0410;
            10'h1F5 : data_reg <= 16'h4C13;
            10'h1F6 : data_reg <= 16'h4E08;
            10'h1F7 : data_reg <= 16'h3CF0;
            10'h1F8 : data_reg <= 16'h3D2B;
            10'h1F9 : data_reg <= 16'h352C;
            10'h1FA : data_reg <= 16'h2D3C;
            10'h1FB : data_reg <= 16'h2C3B;
            10'h1FC : data_reg <= 16'h3D10;
            10'h1FD : data_reg <= 16'h0000;
            10'h1FE : data_reg <= 16'h3C12;
            10'h1FF : data_reg <= 16'h4C12;
            10'h200 : data_reg <= 16'h3E4E;
            10'h201 : data_reg <= 16'h041C;
            10'h202 : data_reg <= 16'h4C13;
            10'h203 : data_reg <= 16'h4E08;
            10'h204 : data_reg <= 16'h3CF0;
            10'h205 : data_reg <= 16'h3D2B;
            10'h206 : data_reg <= 16'h362C;
            10'h207 : data_reg <= 16'h3310;
            10'h208 : data_reg <= 16'hD221;
            10'h209 : data_reg <= 16'h0926;
            10'h20A : data_reg <= 16'h5221;
            10'h20B : data_reg <= 16'h1131;
            10'h20C : data_reg <= 16'h3343;
            10'h20D : data_reg <= 16'h3E25;
            10'h20E : data_reg <= 16'h3221;
            10'h20F : data_reg <= 16'h3123;
            10'h210 : data_reg <= 16'h0A3C;
            10'h211 : data_reg <= 16'h2C36;
            10'h212 : data_reg <= 16'h0A3C;
            10'h213 : data_reg <= 16'h2C35;
            10'h214 : data_reg <= 16'h0A3C;
            10'h215 : data_reg <= 16'h2C33;
            10'h216 : data_reg <= 16'h3C0D;
            10'h217 : data_reg <= 16'h0B23;
            10'h218 : data_reg <= 16'h3C2C;
            10'h219 : data_reg <= 16'h0B24;
            10'h21A : data_reg <= 16'h3C2C;
            10'h21B : data_reg <= 16'h0B25;
            10'h21C : data_reg <= 16'h3C2C;
            10'h21D : data_reg <= 16'h0B26;
            10'h21E : data_reg <= 16'h3C2C;
            10'h21F : data_reg <= 16'h0B27;
            10'h220 : data_reg <= 16'h3C2C;
            10'h221 : data_reg <= 16'h3B2D;
            10'h222 : data_reg <= 16'h102C;
            10'h223 : data_reg <= 16'h003D;
            10'h224 : data_reg <= 16'h0000;
            10'h225 : data_reg <= 16'h3C12;
            10'h226 : data_reg <= 16'h4C12;
            10'h227 : data_reg <= 16'h3E4E;
            10'h228 : data_reg <= 16'h04B3;
            10'h229 : data_reg <= 16'h4C13;
            10'h22A : data_reg <= 16'h4E08;
            10'h22B : data_reg <= 16'h3CF0;
            10'h22C : data_reg <= 16'h3D2B;
            10'h22D : data_reg <= 16'h352C;
            10'h22E : data_reg <= 16'h2D3C;
            10'h22F : data_reg <= 16'h2C3B;
            10'h230 : data_reg <= 16'h3D10;
            10'h231 : data_reg <= 16'h0000;
            10'h232 : data_reg <= 16'h3C12;
            10'h233 : data_reg <= 16'h4C12;
            10'h234 : data_reg <= 16'h3E4E;
            10'h235 : data_reg <= 16'h0494;
            10'h236 : data_reg <= 16'h4C13;
            10'h237 : data_reg <= 16'h4E08;
            10'h238 : data_reg <= 16'h3CF0;
            10'h239 : data_reg <= 16'h3D2B;
            10'h23A : data_reg <= 16'h362C;
            10'h23B : data_reg <= 16'h2D3C;
            10'h23C : data_reg <= 16'h2C3B;
            10'h23D : data_reg <= 16'h3D10;
            10'h23E : data_reg <= 16'h0000;
            10'h23F : data_reg <= 16'h3C12;
            10'h240 : data_reg <= 16'h4C12;
            10'h241 : data_reg <= 16'h3E4E;
            10'h242 : data_reg <= 16'h0367;
            10'h243 : data_reg <= 16'h4C13;
            10'h244 : data_reg <= 16'h4E08;
            10'h245 : data_reg <= 16'h3CF0;
            10'h246 : data_reg <= 16'h3D2B;
            10'h247 : data_reg <= 16'h372C;
            10'h248 : data_reg <= 16'h3311;
            10'h249 : data_reg <= 16'h3410;
            10'h24A : data_reg <= 16'hC224;
            10'h24B : data_reg <= 16'h0925;
            10'h24C : data_reg <= 16'h4411;
            10'h24D : data_reg <= 16'h3C34;
            10'h24E : data_reg <= 16'h0B21;
            10'h24F : data_reg <= 16'h3C2C;
            10'h250 : data_reg <= 16'h0B22;
            10'h251 : data_reg <= 16'h232C;
            10'h252 : data_reg <= 16'h2732;
            10'h253 : data_reg <= 16'h210C;
            10'h254 : data_reg <= 16'h3C33;
            10'h255 : data_reg <= 16'h320A;
            10'h256 : data_reg <= 16'h3C2C;
            10'h257 : data_reg <= 16'h310A;
            10'h258 : data_reg <= 16'h262C;
            10'h259 : data_reg <= 16'h233E;
            10'h25A : data_reg <= 16'h3C31;
            10'h25B : data_reg <= 16'h370A;
            10'h25C : data_reg <= 16'h3C2C;
            10'h25D : data_reg <= 16'h360A;
            10'h25E : data_reg <= 16'h3C2C;
            10'h25F : data_reg <= 16'h350A;
            10'h260 : data_reg <= 16'h3C2C;
            10'h261 : data_reg <= 16'h340A;
            10'h262 : data_reg <= 16'h3C2C;
            10'h263 : data_reg <= 16'h330A;
            10'h264 : data_reg <= 16'h0D2C;
            10'h265 : data_reg <= 16'h223C;
            10'h266 : data_reg <= 16'h2C0B;
            10'h267 : data_reg <= 16'h233C;
            10'h268 : data_reg <= 16'h2C0B;
            10'h269 : data_reg <= 16'h243C;
            10'h26A : data_reg <= 16'h2C0B;
            10'h26B : data_reg <= 16'h253C;
            10'h26C : data_reg <= 16'h2C0B;
            10'h26D : data_reg <= 16'h352D;
            10'h26E : data_reg <= 16'h3D16;
            10'h26F : data_reg <= 16'h3221;
            10'h270 : data_reg <= 16'h2D3C;
            10'h271 : data_reg <= 16'h2C3B;
            10'h272 : data_reg <= 16'h3D10;
            10'h273 : data_reg <= 16'h0000;
            10'h274 : data_reg <= 16'h3C12;
            10'h275 : data_reg <= 16'h4C12;
            10'h276 : data_reg <= 16'h3E4E;
            10'h277 : data_reg <= 16'h04FC;
            10'h278 : data_reg <= 16'h4C13;
            10'h279 : data_reg <= 16'h4E08;
            10'h27A : data_reg <= 16'h3CF0;
            10'h27B : data_reg <= 16'h3D2B;
            10'h27C : data_reg <= 16'h332C;
            10'h27D : data_reg <= 16'h3410;
            10'h27E : data_reg <= 16'hC4F2;
            10'h27F : data_reg <= 16'h1101;
            10'h280 : data_reg <= 16'h3242;
            10'h281 : data_reg <= 16'h0923;
            10'h282 : data_reg <= 16'h3311;
            10'h283 : data_reg <= 16'h5322;
            10'h284 : data_reg <= 16'h3151;
            10'h285 : data_reg <= 16'h3D25;
            10'h286 : data_reg <= 16'h0A3C;
            10'h287 : data_reg <= 16'h2C35;
            10'h288 : data_reg <= 16'h0A3C;
            10'h289 : data_reg <= 16'h2C34;
            10'h28A : data_reg <= 16'h0A3C;
            10'h28B : data_reg <= 16'h2C33;
            10'h28C : data_reg <= 16'h0A3C;
            10'h28D : data_reg <= 16'h2C32;
            10'h28E : data_reg <= 16'h3C0D;
            10'h28F : data_reg <= 16'h0B21;
            10'h290 : data_reg <= 16'h3C2C;
            10'h291 : data_reg <= 16'h0B22;
            10'h292 : data_reg <= 16'h3C2C;
            10'h293 : data_reg <= 16'h0B23;
            10'h294 : data_reg <= 16'h3C2C;
            10'h295 : data_reg <= 16'h0B25;
            10'h296 : data_reg <= 16'h3C2C;
            10'h297 : data_reg <= 16'h0B26;
            10'h298 : data_reg <= 16'h3C2C;
            10'h299 : data_reg <= 16'h0B24;
            10'h29A : data_reg <= 16'h3C2C;
            10'h29B : data_reg <= 16'h342D;
            10'h29C : data_reg <= 16'h162C;
            10'h29D : data_reg <= 16'h3C3D;
            10'h29E : data_reg <= 16'h3B2D;
            10'h29F : data_reg <= 16'h102C;
            10'h2A0 : data_reg <= 16'h003D;
            10'h2A1 : data_reg <= 16'h0000;
            10'h2A2 : data_reg <= 16'h3C12;
            10'h2A3 : data_reg <= 16'h4C12;
            10'h2A4 : data_reg <= 16'h3E4E;
            10'h2A5 : data_reg <= 16'h0572;
            10'h2A6 : data_reg <= 16'h4C13;
            10'h2A7 : data_reg <= 16'h4E08;
            10'h2A8 : data_reg <= 16'h3CF0;
            10'h2A9 : data_reg <= 16'h3D2B;
            10'h2AA : data_reg <= 16'h352C;
            10'h2AB : data_reg <= 16'h2D3C;
            10'h2AC : data_reg <= 16'h2C3B;
            10'h2AD : data_reg <= 16'h3D10;
            10'h2AE : data_reg <= 16'h0000;
            10'h2AF : data_reg <= 16'h3C12;
            10'h2B0 : data_reg <= 16'h4C12;
            10'h2B1 : data_reg <= 16'h3E4E;
            10'h2B2 : data_reg <= 16'h0580;
            10'h2B3 : data_reg <= 16'h4C13;
            10'h2B4 : data_reg <= 16'h4E08;
            10'h2B5 : data_reg <= 16'h3CF0;
            10'h2B6 : data_reg <= 16'h3D2B;
            10'h2B7 : data_reg <= 16'h362C;
            10'h2B8 : data_reg <= 16'h3C11;
            10'h2B9 : data_reg <= 16'hC210;
            10'h2BA : data_reg <= 16'h0926;
            10'h2BB : data_reg <= 16'hE123;
            10'h2BC : data_reg <= 16'h4C21;
            10'h2BD : data_reg <= 16'h2231;
            10'h2BE : data_reg <= 16'h325C;
            10'h2BF : data_reg <= 16'h3E25;
            10'h2C0 : data_reg <= 16'h3D24;
            10'h2C1 : data_reg <= 16'h0A3C;
            10'h2C2 : data_reg <= 16'h2C34;
            10'h2C3 : data_reg <= 16'h0A3C;
            10'h2C4 : data_reg <= 16'h2C36;
            10'h2C5 : data_reg <= 16'h0A3C;
            10'h2C6 : data_reg <= 16'h2C34;
            10'h2C7 : data_reg <= 16'h0A3C;
            10'h2C8 : data_reg <= 16'h2C33;
            10'h2C9 : data_reg <= 16'h0A3C;
            10'h2CA : data_reg <= 16'h2C32;
            10'h2CB : data_reg <= 16'h0A3C;
            10'h2CC : data_reg <= 16'h2C31;
            10'h2CD : data_reg <= 16'h3C0D;
            10'h2CE : data_reg <= 16'h0B22;
            10'h2CF : data_reg <= 16'h3C2C;
            10'h2D0 : data_reg <= 16'h0B23;
            10'h2D1 : data_reg <= 16'h3C2C;
            10'h2D2 : data_reg <= 16'h0B24;
            10'h2D3 : data_reg <= 16'h3C2C;
            10'h2D4 : data_reg <= 16'h0B25;
            10'h2D5 : data_reg <= 16'h3C2C;
            10'h2D6 : data_reg <= 16'h0B26;
            10'h2D7 : data_reg <= 16'h3C2C;
            10'h2D8 : data_reg <= 16'h0B27;
            10'h2D9 : data_reg <= 16'h3C2C;
            10'h2DA : data_reg <= 16'h0B28;
            10'h2DB : data_reg <= 16'h3C2C;
            10'h2DC : data_reg <= 16'h0B21;
            10'h2DD : data_reg <= 16'h3C2C;
            10'h2DE : data_reg <= 16'h3B2D;
            10'h2DF : data_reg <= 16'h102C;
            10'h2E0 : data_reg <= 16'h003D;
            10'h2E1 : data_reg <= 16'h0000;
            10'h2E2 : data_reg <= 16'h3C12;
            10'h2E3 : data_reg <= 16'h4C12;
            10'h2E4 : data_reg <= 16'h3E4E;
            10'h2E5 : data_reg <= 16'h04CA;
            10'h2E6 : data_reg <= 16'h4C13;
            10'h2E7 : data_reg <= 16'h4E08;
            10'h2E8 : data_reg <= 16'h3CF0;
            10'h2E9 : data_reg <= 16'h3D2B;
            10'h2EA : data_reg <= 16'h0C2C;
            10'h2EB : data_reg <= 16'h3221;
            10'h2EC : data_reg <= 16'h0A3C;
            10'h2ED : data_reg <= 16'h2C31;
            10'h2EE : data_reg <= 16'h3310;
            10'h2EF : data_reg <= 16'h3C11;
            10'h2F0 : data_reg <= 16'hBC22;
            10'h2F1 : data_reg <= 16'h3C34;
            10'h2F2 : data_reg <= 16'h3B2D;
            10'h2F3 : data_reg <= 16'h102C;
            10'h2F4 : data_reg <= 16'h003D;
            10'h2F5 : data_reg <= 16'h0000;
            10'h2F6 : data_reg <= 16'h3C12;
            10'h2F7 : data_reg <= 16'h4C12;
            10'h2F8 : data_reg <= 16'h3E4E;
            10'h2F9 : data_reg <= 16'h061E;
            10'h2FA : data_reg <= 16'h4C13;
            10'h2FB : data_reg <= 16'h4E08;
            10'h2FC : data_reg <= 16'h3CF0;
            10'h2FD : data_reg <= 16'h3D2B;
            10'h2FE : data_reg <= 16'h352C;
            10'h2FF : data_reg <= 16'h2D3C;
            10'h300 : data_reg <= 16'h2C3B;
            10'h301 : data_reg <= 16'h3D10;
            10'h302 : data_reg <= 16'h0000;
            10'h303 : data_reg <= 16'h3C12;
            10'h304 : data_reg <= 16'h4C12;
            10'h305 : data_reg <= 16'h3E4E;
            10'h306 : data_reg <= 16'h0639;
            10'h307 : data_reg <= 16'h4C13;
            10'h308 : data_reg <= 16'h4E08;
            10'h309 : data_reg <= 16'h3CF0;
            10'h30A : data_reg <= 16'h3D2B;
            10'h30B : data_reg <= 16'h362C;
            10'h30C : data_reg <= 16'h2D3C;
            10'h30D : data_reg <= 16'h2C37;
            10'h30E : data_reg <= 16'h3D16;
            10'h30F : data_reg <= 16'hC423;
            10'h310 : data_reg <= 16'h0926;
            10'h311 : data_reg <= 16'h4321;
            10'h312 : data_reg <= 16'hF03B;
            10'h313 : data_reg <= 16'h110B;
            10'h314 : data_reg <= 16'h213C;
            10'h315 : data_reg <= 16'h5342;
            10'h316 : data_reg <= 16'h3C5C;
            10'h317 : data_reg <= 16'h38FC;
            10'h318 : data_reg <= 16'hEC0A;
            10'h319 : data_reg <= 16'hEB28;
            10'h31A : data_reg <= 16'h4311;
            10'h31B : data_reg <= 16'h2533;
            10'h31C : data_reg <= 16'h273E;
            10'h31D : data_reg <= 16'h3C3D;
            10'h31E : data_reg <= 16'h380A;
            10'h31F : data_reg <= 16'h3C2C;
            10'h320 : data_reg <= 16'h370A;
            10'h321 : data_reg <= 16'h3C2C;
            10'h322 : data_reg <= 16'h360A;
            10'h323 : data_reg <= 16'h3C2C;
            10'h324 : data_reg <= 16'h350A;
            10'h325 : data_reg <= 16'h3C2C;
            10'h326 : data_reg <= 16'h340A;
            10'h327 : data_reg <= 16'h3C2C;
            10'h328 : data_reg <= 16'h330A;
            10'h329 : data_reg <= 16'h3C2C;
            10'h32A : data_reg <= 16'h320A;
            10'h32B : data_reg <= 16'h0D2C;
            10'h32C : data_reg <= 16'h6548;
            10'h32D : data_reg <= 16'h6C6C;
            10'h32E : data_reg <= 16'h2C6F;
            10'h32F : data_reg <= 16'h7720;
            10'h330 : data_reg <= 16'h726F;
            10'h331 : data_reg <= 16'h646C;
            10'h332 : data_reg <= 16'h0D21;
            10'h333 : data_reg <= 16'h000A;
            10'h334 : data_reg <= 16'h2D3C;
            10'h335 : data_reg <= 16'h2C3B;
            10'h336 : data_reg <= 16'h3D10;
            10'h337 : data_reg <= 16'h0000;
            10'h338 : data_reg <= 16'h3C12;
            10'h339 : data_reg <= 16'h4C12;
            10'h33A : data_reg <= 16'h3E4E;
            10'h33B : data_reg <= 16'h0658;
            10'h33C : data_reg <= 16'h4C13;
            10'h33D : data_reg <= 16'h4E08;
            10'h33E : data_reg <= 16'h3CF0;
            10'h33F : data_reg <= 16'h3D2B;
            10'h340 : data_reg <= 16'h312C;
            10'h341 : data_reg <= 16'h2D3C;
            10'h342 : data_reg <= 16'h2C3B;
            10'h343 : data_reg <= 16'h3D10;
            10'h344 : data_reg <= 16'h0000;
            10'h345 : data_reg <= 16'h3C12;
            10'h346 : data_reg <= 16'h4C12;
            10'h347 : data_reg <= 16'h3E4E;
            10'h348 : data_reg <= 16'h018B;
            10'h349 : data_reg <= 16'h4C13;
            10'h34A : data_reg <= 16'h4E08;
            10'h34B : data_reg <= 16'h3CF0;
            10'h34C : data_reg <= 16'h3D2B;
            10'h34D : data_reg <= 16'h0C2C;
            10'h34E : data_reg <= 16'h000E;
            default : data_reg <= 0;
        endcase
    assign data_out = ( enable ? data_reg : 0 );
endmodule
