`define test_instruction_bin_size 938
`define test_instruction_bin 7504'h00e8e10c1d0b1cd03ee53c23009f1e3e3c22001c221d6d8c9c6d8c221c281b0de10c1d0b1cd03ee53c2301071e3e3c22001c221d6d8c9c6d8c221c281b0de10c1d0b1cd03ee53c2300361e3e3c221c221d6d8c9c6d8c221c281b0d1fd00c1d0b1cd03ee53c23002e1e3e3c22001c221d6d8c9c6d8c221c281b0de2e10a112ae8e2e10a11e7d120c1e70c1d0b1cd03ee53c23ffff1e3e3c22001c221d6d8c9c6d8c221c281b0d113f28e0e60c1d0b1cd03ee53c23032a1e3e3c22001c221d6d8c9c6d8c221c281b0da1211121e10c1d0b1cd03ee53c23032b1e3e3c221c221d6d8c9c6d8c221c281b0de10a11e55c2d1c8c201c24e10a11e320e45c201c8c251c24e10a11df20cf5c2a1c8c251c241e0c1d0b1cd03ee53c23032a1e3e3c22001c221d6d8c9c6d8c221c281b0de00c1d0b1cd03ee53c23029c1e3e3c22001c221d6d8c9c6d8c221c281b0db120e00c1d0b1cd03ee53c23032a1e3e3c22001c221d6d8c9c6d8c221c281b0db121e00c1d0b1cd03ee53c23032a1e3e3c22001c221d6d8c9c6d8c221c281b0da1201e0c1d0b1cd03ee53c23032a1e3e3c22001c221d6d8c9c6d8c221c281b0de00c1d0b1cd03ee53c23021e1e3e3c221c221d6d8c9c6d8c221c281b0da1211121e10a119226e10a1182271221e10a1172e10a11632e132de10a11525c251c8c251c24125c2a1c8c2a1c24e10a114222e10a11425c251c8c251c24125c2a1c8c2a1c24e10a11e532e55c221c8c231c24e10a11e532e55c281c8c2c1c24125c241c8c261c24e10a11315c2f1c8c201c24115c2a1c8c201c24e10a1102120c1d0b1cd03ee53c230c801e3e3c22001c221d6d8c9c6d8c221c281b0de10a11261a0c1d0b1cd03ee53c2300301e3e3c221c221d6d8c9c6d8c221c281b0d19d00c1d0b1cd03ee53c23002a1e3e3c221c221d6d8c9c6d8c221c281b0de2e00c1d0b1cd03ee53c2300dd1e3e3c22001c221d6d8c9c6d8c221c281b0de6a302133321113122e9d1132012d00c1d0b1cd03ee53c23002c1e3e3c221c221d6d8c9c6d8c221c281b0d11d00c1d0b1cd03ee53c23002a1e3e3c221c221d6d8c9c6d8c221c281b0de2e00c1d0b1cd03ee53c2300751e3e3c22001c221d6d8c9c6d8c221c281b0de6a302133321113122c120132012d00c1d0b1cd03ee53c23002c1e3e3c221c221d6d8c9c6d8c221c281b0d11d00c1d0b1cd03ee53c23002a1e3e3c22001c221d6d8c9c6d8c221c281b0de2193922c9019000001480001e0c1d0b1cd03ee53c2303301e3e3c221c221d6d8c9c6d8c221c281b0d1d6d8c9c6d8c221c284d525341
