module rom4(input clk, input enable, input [8-1:0] addr, output [8-1:0] data);
    reg [8-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            8'h0 : data_reg <= 8'h41;
            8'h1 : data_reg <= 8'h53;
            8'h2 : data_reg <= 8'h52;
            8'h3 : data_reg <= 8'h4D;
            8'h4 : data_reg <= 8'h3C;
            8'h5 : data_reg <= 8'h2D;
            8'h6 : data_reg <= 8'h3B;
            8'h7 : data_reg <= 8'h2C;
            8'h8 : data_reg <= 8'h10;
            8'h9 : data_reg <= 8'h3D;
            8'hA : data_reg <= 8'h11;
            8'hB : data_reg <= 8'h3C;
            8'hC : data_reg <= 8'h00;
            8'hD : data_reg <= 8'h00;
            8'hE : data_reg <= 8'h00;
            8'hF : data_reg <= 8'h00;
            8'h10 : data_reg <= 8'h12;
            8'h11 : data_reg <= 8'h4C;
            8'h12 : data_reg <= 8'h4E;
            8'h13 : data_reg <= 8'h3E;
            8'h14 : data_reg <= 8'h9A;
            8'h15 : data_reg <= 8'h13;
            8'h16 : data_reg <= 8'h4C;
            8'h17 : data_reg <= 8'h08;
            8'h18 : data_reg <= 8'h4E;
            8'h19 : data_reg <= 8'hF0;
            8'h1A : data_reg <= 8'h3C;
            8'h1B : data_reg <= 8'h2B;
            8'h1C : data_reg <= 8'h3D;
            8'h1D : data_reg <= 8'h2C;
            8'h1E : data_reg <= 8'h3F;
            8'h1F : data_reg <= 8'h3C;
            8'h20 : data_reg <= 8'h2D;
            8'h21 : data_reg <= 8'h3B;
            8'h22 : data_reg <= 8'h2C;
            8'h23 : data_reg <= 8'h10;
            8'h24 : data_reg <= 8'h3D;
            8'h25 : data_reg <= 8'h11;
            8'h26 : data_reg <= 8'h3C;
            8'h27 : data_reg <= 8'h00;
            8'h28 : data_reg <= 8'h00;
            8'h29 : data_reg <= 8'h00;
            8'h2A : data_reg <= 8'h00;
            8'h2B : data_reg <= 8'h12;
            8'h2C : data_reg <= 8'h4C;
            8'h2D : data_reg <= 8'h4E;
            8'h2E : data_reg <= 8'h3E;
            8'h2F : data_reg <= 8'h4E;
            8'h30 : data_reg <= 8'h13;
            8'h31 : data_reg <= 8'h4C;
            8'h32 : data_reg <= 8'h08;
            8'h33 : data_reg <= 8'h4E;
            8'h34 : data_reg <= 8'hF0;
            8'h35 : data_reg <= 8'h3C;
            8'h36 : data_reg <= 8'h2B;
            8'h37 : data_reg <= 8'h3D;
            8'h38 : data_reg <= 8'h2C;
            8'h39 : data_reg <= 8'h3E;
            8'h3A : data_reg <= 8'h34;
            8'h3B : data_reg <= 8'h13;
            8'h3C : data_reg <= 8'h42;
            8'h3D : data_reg <= 8'h35;
            8'h3E : data_reg <= 8'hF5;
            8'h3F : data_reg <= 8'h33;
            8'h40 : data_reg <= 8'h11;
            8'h41 : data_reg <= 8'h42;
            8'h42 : data_reg <= 8'h35;
            8'h43 : data_reg <= 8'h23;
            8'h44 : data_reg <= 8'hE5;
            8'h45 : data_reg <= 8'h10;
            8'h46 : data_reg <= 8'hE2;
            8'h47 : data_reg <= 8'h13;
            8'h48 : data_reg <= 8'h41;
            8'h49 : data_reg <= 8'h33;
            8'h4A : data_reg <= 8'h10;
            8'h4B : data_reg <= 8'hE3;
            8'h4C : data_reg <= 8'h24;
            8'h4D : data_reg <= 8'h02;
            8'h4E : data_reg <= 8'h14;
            8'h4F : data_reg <= 8'h3C;
            8'h50 : data_reg <= 8'h1E;
            8'h51 : data_reg <= 8'hAC;
            8'h52 : data_reg <= 8'h3C;
            8'h53 : data_reg <= 8'h1D;
            8'h54 : data_reg <= 8'h7C;
            8'h55 : data_reg <= 8'h31;
            8'h56 : data_reg <= 8'h12;
            8'h57 : data_reg <= 8'hE1;
            8'h58 : data_reg <= 8'h3C;
            8'h59 : data_reg <= 8'h2D;
            8'h5A : data_reg <= 8'h3B;
            8'h5B : data_reg <= 8'h2C;
            8'h5C : data_reg <= 8'h10;
            8'h5D : data_reg <= 8'h3D;
            8'h5E : data_reg <= 8'h11;
            8'h5F : data_reg <= 8'h3C;
            8'h60 : data_reg <= 8'h00;
            8'h61 : data_reg <= 8'h00;
            8'h62 : data_reg <= 8'h00;
            8'h63 : data_reg <= 8'h00;
            8'h64 : data_reg <= 8'h12;
            8'h65 : data_reg <= 8'h4C;
            8'h66 : data_reg <= 8'h4E;
            8'h67 : data_reg <= 8'h3E;
            8'h68 : data_reg <= 8'h3A;
            8'h69 : data_reg <= 8'h13;
            8'h6A : data_reg <= 8'h4C;
            8'h6B : data_reg <= 8'h08;
            8'h6C : data_reg <= 8'h4E;
            8'h6D : data_reg <= 8'hF0;
            8'h6E : data_reg <= 8'h3C;
            8'h6F : data_reg <= 8'h2B;
            8'h70 : data_reg <= 8'h3D;
            8'h71 : data_reg <= 8'h2C;
            8'h72 : data_reg <= 8'h04;
            8'h73 : data_reg <= 8'h18;
            8'h74 : data_reg <= 8'h3D;
            8'h75 : data_reg <= 8'h14;
            8'h76 : data_reg <= 8'h3C;
            8'h77 : data_reg <= 8'h1F;
            8'h78 : data_reg <= 8'hAC;
            8'h79 : data_reg <= 8'h3C;
            8'h7A : data_reg <= 8'h1C;
            8'h7B : data_reg <= 8'h7C;
            8'h7C : data_reg <= 8'h32;
            8'h7D : data_reg <= 8'h3C;
            8'h7E : data_reg <= 8'h2D;
            8'h7F : data_reg <= 8'h3B;
            8'h80 : data_reg <= 8'h2C;
            8'h81 : data_reg <= 8'h10;
            8'h82 : data_reg <= 8'h3D;
            8'h83 : data_reg <= 8'h11;
            8'h84 : data_reg <= 8'h3C;
            8'h85 : data_reg <= 8'h00;
            8'h86 : data_reg <= 8'h00;
            8'h87 : data_reg <= 8'h00;
            8'h88 : data_reg <= 8'h00;
            8'h89 : data_reg <= 8'h12;
            8'h8A : data_reg <= 8'h4C;
            8'h8B : data_reg <= 8'h4E;
            8'h8C : data_reg <= 8'h3E;
            8'h8D : data_reg <= 8'h97;
            8'h8E : data_reg <= 8'h13;
            8'h8F : data_reg <= 8'h4C;
            8'h90 : data_reg <= 8'h08;
            8'h91 : data_reg <= 8'h4E;
            8'h92 : data_reg <= 8'hF0;
            8'h93 : data_reg <= 8'h3C;
            8'h94 : data_reg <= 8'h2B;
            8'h95 : data_reg <= 8'h3D;
            8'h96 : data_reg <= 8'h2C;
            8'h97 : data_reg <= 8'h00;
            8'h98 : data_reg <= 8'h00;
            8'h99 : data_reg <= 8'h3E;
            default : data_reg <= 0;
        endcase
    assign data = ( enable ? data_reg : 0 );
endmodule
