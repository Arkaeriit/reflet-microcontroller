../submodules/reflet/rtl/reflet.vh