//The code used to make this ROM is in software/helloWorld.asm
module rom2(input clk, input enable ,input [10:0] addr, output [7:0] data_out);
reg [7:0] ret; assign data_out = (enable ? ret : 8'h0);
always @ (posedge clk)
case(addr)
  11'h0 : ret <= 8'h41;
  11'h1 : ret <= 8'h53;
  11'h2 : ret <= 8'h52;
  11'h3 : ret <= 8'h4d;
  11'h4 : ret <= 8'h14;
  11'h5 : ret <= 8'h3c;
  11'h6 : ret <= 8'h10;
  11'h7 : ret <= 8'h3b;
  11'h8 : ret <= 8'h10;
  11'h9 : ret <= 8'h7b;
  11'ha : ret <= 8'hac;
  11'hb : ret <= 8'h3b;
  11'hc : ret <= 8'h14;
  11'hd : ret <= 8'h7b;
  11'he : ret <= 8'hac;
  11'hf : ret <= 8'h3b;
  11'h10 : ret <= 8'h1b;
  11'h11 : ret <= 8'h7b;
  11'h12 : ret <= 8'hac;
  11'h13 : ret <= 8'h3b;
  11'h14 : ret <= 8'h15;
  11'h15 : ret <= 8'h7b;
  11'h16 : ret <= 8'h3f;
  11'h17 : ret <= 8'h14;
  11'h18 : ret <= 8'h3c;
  11'h19 : ret <= 8'h10;
  11'h1a : ret <= 8'h3b;
  11'h1b : ret <= 8'h10;
  11'h1c : ret <= 8'h7b;
  11'h1d : ret <= 8'hac;
  11'h1e : ret <= 8'h3b;
  11'h1f : ret <= 8'h10;
  11'h20 : ret <= 8'h7b;
  11'h21 : ret <= 8'hac;
  11'h22 : ret <= 8'h3b;
  11'h23 : ret <= 8'h13;
  11'h24 : ret <= 8'h7b;
  11'h25 : ret <= 8'hac;
  11'h26 : ret <= 8'h3b;
  11'h27 : ret <= 8'h1a;
  11'h28 : ret <= 8'h7b;
  11'h29 : ret <= 8'h8;
  11'h2a : ret <= 8'h48;
  11'h2b : ret <= 8'h65;
  11'h2c : ret <= 8'h6c;
  11'h2d : ret <= 8'h6c;
  11'h2e : ret <= 8'h6f;
  11'h2f : ret <= 8'h2c;
  11'h30 : ret <= 8'h20;
  11'h31 : ret <= 8'h77;
  11'h32 : ret <= 8'h6f;
  11'h33 : ret <= 8'h72;
  11'h34 : ret <= 8'h6c;
  11'h35 : ret <= 8'h64;
  11'h36 : ret <= 8'h21;
  11'h37 : ret <= 8'hd;
  11'h38 : ret <= 8'ha;
  11'h39 : ret <= 8'h0;
  11'h3a : ret <= 8'h14;
  11'h3b : ret <= 8'h3c;
  11'h3c : ret <= 8'h10;
  11'h3d : ret <= 8'h3b;
  11'h3e : ret <= 8'h10;
  11'h3f : ret <= 8'h7b;
  11'h40 : ret <= 8'hac;
  11'h41 : ret <= 8'h3b;
  11'h42 : ret <= 8'h10;
  11'h43 : ret <= 8'h7b;
  11'h44 : ret <= 8'hac;
  11'h45 : ret <= 8'h3b;
  11'h46 : ret <= 8'h17;
  11'h47 : ret <= 8'h7b;
  11'h48 : ret <= 8'hac;
  11'h49 : ret <= 8'h3b;
  11'h4a : ret <= 8'h15;
  11'h4b : ret <= 8'h7b;
  11'h4c : ret <= 8'hf0;
  11'h4d : ret <= 8'h3f;
  11'h4e : ret <= 8'h14;
  11'h4f : ret <= 8'h3c;
  11'h50 : ret <= 8'h10;
  11'h51 : ret <= 8'h3b;
  11'h52 : ret <= 8'h10;
  11'h53 : ret <= 8'h7b;
  11'h54 : ret <= 8'hac;
  11'h55 : ret <= 8'h3b;
  11'h56 : ret <= 8'h10;
  11'h57 : ret <= 8'h7b;
  11'h58 : ret <= 8'hac;
  11'h59 : ret <= 8'h3b;
  11'h5a : ret <= 8'h12;
  11'h5b : ret <= 8'h7b;
  11'h5c : ret <= 8'hac;
  11'h5d : ret <= 8'h3b;
  11'h5e : ret <= 8'h1a;
  11'h5f : ret <= 8'h7b;
  11'h60 : ret <= 8'h31;
  11'h61 : ret <= 8'h14;
  11'h62 : ret <= 8'h3c;
  11'h63 : ret <= 8'h10;
  11'h64 : ret <= 8'h3b;
  11'h65 : ret <= 8'h10;
  11'h66 : ret <= 8'h7b;
  11'h67 : ret <= 8'hac;
  11'h68 : ret <= 8'h3b;
  11'h69 : ret <= 8'h13;
  11'h6a : ret <= 8'h7b;
  11'h6b : ret <= 8'hac;
  11'h6c : ret <= 8'h3b;
  11'h6d : ret <= 8'h17;
  11'h6e : ret <= 8'h7b;
  11'h6f : ret <= 8'hac;
  11'h70 : ret <= 8'h3b;
  11'h71 : ret <= 8'h11;
  11'h72 : ret <= 8'h7b;
  11'h73 : ret <= 8'hc;
  11'h74 : ret <= 8'he;
  11'h75 : ret <= 8'h0;
  11'h76 : ret <= 8'h80;
  11'h77 : ret <= 8'h0;
  11'h78 : ret <= 8'hff;
  11'h79 : ret <= 8'h4;
  11'h7a : ret <= 8'hff;
  11'h7b : ret <= 8'h8;
  11'h7c : ret <= 8'hff;
  11'h7d : ret <= 8'h10;
  11'h7e : ret <= 8'hff;
  11'h7f : ret <= 8'h13;
  11'h80 : ret <= 8'hff;
  11'h81 : ret <= 8'h16;
  11'h82 : ret <= 8'hff;
  11'h83 : ret <= 8'h1a;
  11'h84 : ret <= 8'hff;
  11'h85 : ret <= 8'h1c;
  11'h86 : ret <= 8'hff;
  11'h87 : ret <= 8'h22;
  11'h88 : ret <= 8'hb;
  11'h89 : ret <= 8'h24;
  11'h8a : ret <= 8'hb;
  11'h8b : ret <= 8'h14;
  11'h8c : ret <= 8'h3c;
  11'h8d : ret <= 8'h10;
  11'h8e : ret <= 8'h3b;
  11'h8f : ret <= 8'h10;
  11'h90 : ret <= 8'h7b;
  11'h91 : ret <= 8'hac;
  11'h92 : ret <= 8'h3b;
  11'h93 : ret <= 8'h10;
  11'h94 : ret <= 8'h7b;
  11'h95 : ret <= 8'hac;
  11'h96 : ret <= 8'h3b;
  11'h97 : ret <= 8'h18;
  11'h98 : ret <= 8'h7b;
  11'h99 : ret <= 8'hac;
  11'h9a : ret <= 8'h3b;
  11'h9b : ret <= 8'h11;
  11'h9c : ret <= 8'h7b;
  11'h9d : ret <= 8'hf0;
  11'h9e : ret <= 8'h32;
  11'h9f : ret <= 8'h14;
  11'ha0 : ret <= 8'h3c;
  11'ha1 : ret <= 8'h10;
  11'ha2 : ret <= 8'h3b;
  11'ha3 : ret <= 8'h10;
  11'ha4 : ret <= 8'h7b;
  11'ha5 : ret <= 8'hac;
  11'ha6 : ret <= 8'h3b;
  11'ha7 : ret <= 8'h10;
  11'ha8 : ret <= 8'h7b;
  11'ha9 : ret <= 8'hac;
  11'haa : ret <= 8'h3b;
  11'hab : ret <= 8'h1b;
  11'hac : ret <= 8'h7b;
  11'had : ret <= 8'hac;
  11'hae : ret <= 8'h3b;
  11'haf : ret <= 8'h12;
  11'hb0 : ret <= 8'h7b;
  11'hb1 : ret <= 8'h34;
  11'hb2 : ret <= 8'hf2;
  11'hb3 : ret <= 8'h3c;
  11'hb4 : ret <= 8'h10;
  11'hb5 : ret <= 8'hcc;
  11'hb6 : ret <= 8'h24;
  11'hb7 : ret <= 8'h9;
  11'hb8 : ret <= 8'h11;
  11'hb9 : ret <= 8'h42;
  11'hba : ret <= 8'h3c;
  11'hbb : ret <= 8'h21;
  11'hbc : ret <= 8'hec;
  11'hbd : ret <= 8'h10;
  11'hbe : ret <= 8'he2;
  11'hbf : ret <= 8'ha;
  11'hc0 : ret <= 8'h34;
  11'hc1 : ret <= 8'ha;
  11'hc2 : ret <= 8'h32;
  11'hc3 : ret <= 8'hd;
  11'hc4 : ret <= 8'h21;
  11'hc5 : ret <= 8'hb;
  11'hc6 : ret <= 8'h1a;
  11'hc7 : ret <= 8'h31;
  11'hc8 : ret <= 8'h14;
  11'hc9 : ret <= 8'h3c;
  11'hca : ret <= 8'h10;
  11'hcb : ret <= 8'h3b;
  11'hcc : ret <= 8'h10;
  11'hcd : ret <= 8'h7b;
  11'hce : ret <= 8'hac;
  11'hcf : ret <= 8'h3b;
  11'hd0 : ret <= 8'h10;
  11'hd1 : ret <= 8'h7b;
  11'hd2 : ret <= 8'hac;
  11'hd3 : ret <= 8'h3b;
  11'hd4 : ret <= 8'h18;
  11'hd5 : ret <= 8'h7b;
  11'hd6 : ret <= 8'hac;
  11'hd7 : ret <= 8'h3b;
  11'hd8 : ret <= 8'h17;
  11'hd9 : ret <= 8'h7b;
  11'hda : ret <= 8'hc;
  11'hdb : ret <= 8'h1d;
  11'hdc : ret <= 8'h31;
  11'hdd : ret <= 8'h14;
  11'hde : ret <= 8'h3c;
  11'hdf : ret <= 8'h10;
  11'he0 : ret <= 8'h3b;
  11'he1 : ret <= 8'h10;
  11'he2 : ret <= 8'h7b;
  11'he3 : ret <= 8'hac;
  11'he4 : ret <= 8'h3b;
  11'he5 : ret <= 8'h10;
  11'he6 : ret <= 8'h7b;
  11'he7 : ret <= 8'hac;
  11'he8 : ret <= 8'h3b;
  11'he9 : ret <= 8'h18;
  11'hea : ret <= 8'h7b;
  11'heb : ret <= 8'hac;
  11'hec : ret <= 8'h3b;
  11'hed : ret <= 8'h17;
  11'hee : ret <= 8'h7b;
  11'hef : ret <= 8'hc;
  11'hf0 : ret <= 8'ha;
  11'hf1 : ret <= 8'h31;
  11'hf2 : ret <= 8'hd;
  11'hf3 : ret <= 8'h23;
  11'hf4 : ret <= 8'hb;
  11'hf5 : ret <= 8'h24;
  11'hf6 : ret <= 8'hb;
  11'hf7 : ret <= 8'h25;
  11'hf8 : ret <= 8'hb;
  11'hf9 : ret <= 8'h26;
  11'hfa : ret <= 8'hb;
  11'hfb : ret <= 8'h10;
  11'hfc : ret <= 8'h33;
  11'hfd : ret <= 8'h34;
  11'hfe : ret <= 8'h14;
  11'hff : ret <= 8'h3c;
  11'h100 : ret <= 8'h10;
  11'h101 : ret <= 8'h3b;
  11'h102 : ret <= 8'h10;
  11'h103 : ret <= 8'h7b;
  11'h104 : ret <= 8'hac;
  11'h105 : ret <= 8'h3b;
  11'h106 : ret <= 8'h11;
  11'h107 : ret <= 8'h7b;
  11'h108 : ret <= 8'hac;
  11'h109 : ret <= 8'h3b;
  11'h10a : ret <= 8'h13;
  11'h10b : ret <= 8'h7b;
  11'h10c : ret <= 8'hac;
  11'h10d : ret <= 8'h3b;
  11'h10e : ret <= 8'h11;
  11'h10f : ret <= 8'h7b;
  11'h110 : ret <= 8'h35;
  11'h111 : ret <= 8'h14;
  11'h112 : ret <= 8'h3c;
  11'h113 : ret <= 8'h10;
  11'h114 : ret <= 8'h3b;
  11'h115 : ret <= 8'h10;
  11'h116 : ret <= 8'h7b;
  11'h117 : ret <= 8'hac;
  11'h118 : ret <= 8'h3b;
  11'h119 : ret <= 8'h11;
  11'h11a : ret <= 8'h7b;
  11'h11b : ret <= 8'hac;
  11'h11c : ret <= 8'h3b;
  11'h11d : ret <= 8'h12;
  11'h11e : ret <= 8'h7b;
  11'h11f : ret <= 8'hac;
  11'h120 : ret <= 8'h3b;
  11'h121 : ret <= 8'h15;
  11'h122 : ret <= 8'h7b;
  11'h123 : ret <= 8'h36;
  11'h124 : ret <= 8'h10;
  11'h125 : ret <= 8'h24;
  11'h126 : ret <= 8'hc2;
  11'h127 : ret <= 8'h25;
  11'h128 : ret <= 8'h9;
  11'h129 : ret <= 8'h11;
  11'h12a : ret <= 8'h44;
  11'h12b : ret <= 8'h34;
  11'h12c : ret <= 8'h21;
  11'h12d : ret <= 8'h43;
  11'h12e : ret <= 8'h33;
  11'h12f : ret <= 8'h26;
  11'h130 : ret <= 8'h8;
  11'h131 : ret <= 8'h23;
  11'h132 : ret <= 8'h31;
  11'h133 : ret <= 8'ha;
  11'h134 : ret <= 8'h36;
  11'h135 : ret <= 8'ha;
  11'h136 : ret <= 8'h35;
  11'h137 : ret <= 8'ha;
  11'h138 : ret <= 8'h34;
  11'h139 : ret <= 8'ha;
  11'h13a : ret <= 8'h33;
  11'h13b : ret <= 8'hd;
  11'h13c : ret <= 8'h23;
  11'h13d : ret <= 8'hb;
  11'h13e : ret <= 8'h25;
  11'h13f : ret <= 8'hb;
  11'h140 : ret <= 8'h26;
  11'h141 : ret <= 8'hb;
  11'h142 : ret <= 8'h14;
  11'h143 : ret <= 8'h3c;
  11'h144 : ret <= 8'h10;
  11'h145 : ret <= 8'h3b;
  11'h146 : ret <= 8'h10;
  11'h147 : ret <= 8'h7b;
  11'h148 : ret <= 8'hac;
  11'h149 : ret <= 8'h3b;
  11'h14a : ret <= 8'h11;
  11'h14b : ret <= 8'h7b;
  11'h14c : ret <= 8'hac;
  11'h14d : ret <= 8'h3b;
  11'h14e : ret <= 8'h16;
  11'h14f : ret <= 8'h7b;
  11'h150 : ret <= 8'hac;
  11'h151 : ret <= 8'h3b;
  11'h152 : ret <= 8'h1a;
  11'h153 : ret <= 8'h7b;
  11'h154 : ret <= 8'h35;
  11'h155 : ret <= 8'h14;
  11'h156 : ret <= 8'h3c;
  11'h157 : ret <= 8'h10;
  11'h158 : ret <= 8'h3b;
  11'h159 : ret <= 8'h10;
  11'h15a : ret <= 8'h7b;
  11'h15b : ret <= 8'hac;
  11'h15c : ret <= 8'h3b;
  11'h15d : ret <= 8'h11;
  11'h15e : ret <= 8'h7b;
  11'h15f : ret <= 8'hac;
  11'h160 : ret <= 8'h3b;
  11'h161 : ret <= 8'h17;
  11'h162 : ret <= 8'h7b;
  11'h163 : ret <= 8'hac;
  11'h164 : ret <= 8'h3b;
  11'h165 : ret <= 8'h16;
  11'h166 : ret <= 8'h7b;
  11'h167 : ret <= 8'h36;
  11'h168 : ret <= 8'h10;
  11'h169 : ret <= 8'h33;
  11'h16a : ret <= 8'h21;
  11'h16b : ret <= 8'hd2;
  11'h16c : ret <= 8'h26;
  11'h16d : ret <= 8'h9;
  11'h16e : ret <= 8'h21;
  11'h16f : ret <= 8'h52;
  11'h170 : ret <= 8'h31;
  11'h171 : ret <= 8'h11;
  11'h172 : ret <= 8'h43;
  11'h173 : ret <= 8'h33;
  11'h174 : ret <= 8'h25;
  11'h175 : ret <= 8'h8;
  11'h176 : ret <= 8'h21;
  11'h177 : ret <= 8'h32;
  11'h178 : ret <= 8'h23;
  11'h179 : ret <= 8'h31;
  11'h17a : ret <= 8'ha;
  11'h17b : ret <= 8'h36;
  11'h17c : ret <= 8'ha;
  11'h17d : ret <= 8'h35;
  11'h17e : ret <= 8'ha;
  11'h17f : ret <= 8'h33;
  11'h180 : ret <= 8'hd;
  11'h181 : ret <= 8'h23;
  11'h182 : ret <= 8'hb;
  11'h183 : ret <= 8'h24;
  11'h184 : ret <= 8'hb;
  11'h185 : ret <= 8'h25;
  11'h186 : ret <= 8'hb;
  11'h187 : ret <= 8'h26;
  11'h188 : ret <= 8'hb;
  11'h189 : ret <= 8'h27;
  11'h18a : ret <= 8'hb;
  11'h18b : ret <= 8'h14;
  11'h18c : ret <= 8'h3c;
  11'h18d : ret <= 8'h10;
  11'h18e : ret <= 8'h3b;
  11'h18f : ret <= 8'h10;
  11'h190 : ret <= 8'h7b;
  11'h191 : ret <= 8'hac;
  11'h192 : ret <= 8'h3b;
  11'h193 : ret <= 8'h11;
  11'h194 : ret <= 8'h7b;
  11'h195 : ret <= 8'hac;
  11'h196 : ret <= 8'h3b;
  11'h197 : ret <= 8'h1d;
  11'h198 : ret <= 8'h7b;
  11'h199 : ret <= 8'hac;
  11'h19a : ret <= 8'h3b;
  11'h19b : ret <= 8'h1f;
  11'h19c : ret <= 8'h7b;
  11'h19d : ret <= 8'h35;
  11'h19e : ret <= 8'h14;
  11'h19f : ret <= 8'h3c;
  11'h1a0 : ret <= 8'h10;
  11'h1a1 : ret <= 8'h3b;
  11'h1a2 : ret <= 8'h10;
  11'h1a3 : ret <= 8'h7b;
  11'h1a4 : ret <= 8'hac;
  11'h1a5 : ret <= 8'h3b;
  11'h1a6 : ret <= 8'h11;
  11'h1a7 : ret <= 8'h7b;
  11'h1a8 : ret <= 8'hac;
  11'h1a9 : ret <= 8'h3b;
  11'h1aa : ret <= 8'h1c;
  11'h1ab : ret <= 8'h7b;
  11'h1ac : ret <= 8'hac;
  11'h1ad : ret <= 8'h3b;
  11'h1ae : ret <= 8'h18;
  11'h1af : ret <= 8'h7b;
  11'h1b0 : ret <= 8'h36;
  11'h1b1 : ret <= 8'h14;
  11'h1b2 : ret <= 8'h3c;
  11'h1b3 : ret <= 8'h10;
  11'h1b4 : ret <= 8'h3b;
  11'h1b5 : ret <= 8'h10;
  11'h1b6 : ret <= 8'h7b;
  11'h1b7 : ret <= 8'hac;
  11'h1b8 : ret <= 8'h3b;
  11'h1b9 : ret <= 8'h10;
  11'h1ba : ret <= 8'h7b;
  11'h1bb : ret <= 8'hac;
  11'h1bc : ret <= 8'h3b;
  11'h1bd : ret <= 8'h1f;
  11'h1be : ret <= 8'h7b;
  11'h1bf : ret <= 8'hac;
  11'h1c0 : ret <= 8'h3b;
  11'h1c1 : ret <= 8'h13;
  11'h1c2 : ret <= 8'h7b;
  11'h1c3 : ret <= 8'h37;
  11'h1c4 : ret <= 8'h11;
  11'h1c5 : ret <= 8'h33;
  11'h1c6 : ret <= 8'h10;
  11'h1c7 : ret <= 8'h34;
  11'h1c8 : ret <= 8'h24;
  11'h1c9 : ret <= 8'hc2;
  11'h1ca : ret <= 8'h25;
  11'h1cb : ret <= 8'h9;
  11'h1cc : ret <= 8'h11;
  11'h1cd : ret <= 8'h44;
  11'h1ce : ret <= 8'h34;
  11'h1cf : ret <= 8'h21;
  11'h1d0 : ret <= 8'hb;
  11'h1d1 : ret <= 8'h22;
  11'h1d2 : ret <= 8'hb;
  11'h1d3 : ret <= 8'h23;
  11'h1d4 : ret <= 8'h32;
  11'h1d5 : ret <= 8'h27;
  11'h1d6 : ret <= 8'hc;
  11'h1d7 : ret <= 8'h21;
  11'h1d8 : ret <= 8'h33;
  11'h1d9 : ret <= 8'ha;
  11'h1da : ret <= 8'h32;
  11'h1db : ret <= 8'ha;
  11'h1dc : ret <= 8'h31;
  11'h1dd : ret <= 8'h26;
  11'h1de : ret <= 8'h8;
  11'h1df : ret <= 8'h23;
  11'h1e0 : ret <= 8'h31;
  11'h1e1 : ret <= 8'ha;
  11'h1e2 : ret <= 8'h37;
  11'h1e3 : ret <= 8'ha;
  11'h1e4 : ret <= 8'h36;
  11'h1e5 : ret <= 8'ha;
  11'h1e6 : ret <= 8'h35;
  11'h1e7 : ret <= 8'ha;
  11'h1e8 : ret <= 8'h34;
  11'h1e9 : ret <= 8'ha;
  11'h1ea : ret <= 8'h33;
  11'h1eb : ret <= 8'hd;
  11'h1ec : ret <= 8'h22;
  11'h1ed : ret <= 8'hb;
  11'h1ee : ret <= 8'h23;
  11'h1ef : ret <= 8'hb;
  11'h1f0 : ret <= 8'h24;
  11'h1f1 : ret <= 8'hb;
  11'h1f2 : ret <= 8'h25;
  11'h1f3 : ret <= 8'hb;
  11'h1f4 : ret <= 8'h2d;
  11'h1f5 : ret <= 8'h35;
  11'h1f6 : ret <= 8'h16;
  11'h1f7 : ret <= 8'h3d;
  11'h1f8 : ret <= 8'h21;
  11'h1f9 : ret <= 8'h32;
  11'h1fa : ret <= 8'h14;
  11'h1fb : ret <= 8'h3c;
  11'h1fc : ret <= 8'h10;
  11'h1fd : ret <= 8'h3b;
  11'h1fe : ret <= 8'h10;
  11'h1ff : ret <= 8'h7b;
  11'h200 : ret <= 8'hac;
  11'h201 : ret <= 8'h3b;
  11'h202 : ret <= 8'h12;
  11'h203 : ret <= 8'h7b;
  11'h204 : ret <= 8'hac;
  11'h205 : ret <= 8'h3b;
  11'h206 : ret <= 8'h10;
  11'h207 : ret <= 8'h7b;
  11'h208 : ret <= 8'hac;
  11'h209 : ret <= 8'h3b;
  11'h20a : ret <= 8'h1f;
  11'h20b : ret <= 8'h7b;
  11'h20c : ret <= 8'h33;
  11'h20d : ret <= 8'h10;
  11'h20e : ret <= 8'h34;
  11'h20f : ret <= 8'hf2;
  11'h210 : ret <= 8'hc4;
  11'h211 : ret <= 8'h1;
  11'h212 : ret <= 8'h11;
  11'h213 : ret <= 8'h42;
  11'h214 : ret <= 8'h32;
  11'h215 : ret <= 8'h23;
  11'h216 : ret <= 8'h9;
  11'h217 : ret <= 8'h11;
  11'h218 : ret <= 8'h33;
  11'h219 : ret <= 8'h22;
  11'h21a : ret <= 8'h53;
  11'h21b : ret <= 8'h51;
  11'h21c : ret <= 8'h31;
  11'h21d : ret <= 8'h25;
  11'h21e : ret <= 8'h3d;
  11'h21f : ret <= 8'ha;
  11'h220 : ret <= 8'h35;
  11'h221 : ret <= 8'ha;
  11'h222 : ret <= 8'h34;
  11'h223 : ret <= 8'ha;
  11'h224 : ret <= 8'h33;
  11'h225 : ret <= 8'ha;
  11'h226 : ret <= 8'h32;
  11'h227 : ret <= 8'hd;
  11'h228 : ret <= 8'h21;
  11'h229 : ret <= 8'hb;
  11'h22a : ret <= 8'h22;
  11'h22b : ret <= 8'hb;
  11'h22c : ret <= 8'h23;
  11'h22d : ret <= 8'hb;
  11'h22e : ret <= 8'h25;
  11'h22f : ret <= 8'hb;
  11'h230 : ret <= 8'h26;
  11'h231 : ret <= 8'hb;
  11'h232 : ret <= 8'h24;
  11'h233 : ret <= 8'hb;
  11'h234 : ret <= 8'hb;
  11'h235 : ret <= 8'h2d;
  11'h236 : ret <= 8'h34;
  11'h237 : ret <= 8'ha;
  11'h238 : ret <= 8'h16;
  11'h239 : ret <= 8'h3d;
  11'h23a : ret <= 8'h14;
  11'h23b : ret <= 8'h3c;
  11'h23c : ret <= 8'h10;
  11'h23d : ret <= 8'h3b;
  11'h23e : ret <= 8'h10;
  11'h23f : ret <= 8'h7b;
  11'h240 : ret <= 8'hac;
  11'h241 : ret <= 8'h3b;
  11'h242 : ret <= 8'h12;
  11'h243 : ret <= 8'h7b;
  11'h244 : ret <= 8'hac;
  11'h245 : ret <= 8'h3b;
  11'h246 : ret <= 8'h16;
  11'h247 : ret <= 8'h7b;
  11'h248 : ret <= 8'hac;
  11'h249 : ret <= 8'h3b;
  11'h24a : ret <= 8'h12;
  11'h24b : ret <= 8'h7b;
  11'h24c : ret <= 8'h35;
  11'h24d : ret <= 8'h14;
  11'h24e : ret <= 8'h3c;
  11'h24f : ret <= 8'h10;
  11'h250 : ret <= 8'h3b;
  11'h251 : ret <= 8'h10;
  11'h252 : ret <= 8'h7b;
  11'h253 : ret <= 8'hac;
  11'h254 : ret <= 8'h3b;
  11'h255 : ret <= 8'h12;
  11'h256 : ret <= 8'h7b;
  11'h257 : ret <= 8'hac;
  11'h258 : ret <= 8'h3b;
  11'h259 : ret <= 8'h17;
  11'h25a : ret <= 8'h7b;
  11'h25b : ret <= 8'hac;
  11'h25c : ret <= 8'h3b;
  11'h25d : ret <= 8'h10;
  11'h25e : ret <= 8'h7b;
  11'h25f : ret <= 8'h36;
  11'h260 : ret <= 8'h11;
  11'h261 : ret <= 8'h3c;
  11'h262 : ret <= 8'h10;
  11'h263 : ret <= 8'hc2;
  11'h264 : ret <= 8'h26;
  11'h265 : ret <= 8'h9;
  11'h266 : ret <= 8'h23;
  11'h267 : ret <= 8'he1;
  11'h268 : ret <= 8'h21;
  11'h269 : ret <= 8'h4c;
  11'h26a : ret <= 8'h31;
  11'h26b : ret <= 8'h22;
  11'h26c : ret <= 8'h5c;
  11'h26d : ret <= 8'h32;
  11'h26e : ret <= 8'h25;
  11'h26f : ret <= 8'h8;
  11'h270 : ret <= 8'h24;
  11'h271 : ret <= 8'h3d;
  11'h272 : ret <= 8'ha;
  11'h273 : ret <= 8'h34;
  11'h274 : ret <= 8'ha;
  11'h275 : ret <= 8'h36;
  11'h276 : ret <= 8'ha;
  11'h277 : ret <= 8'h34;
  11'h278 : ret <= 8'ha;
  11'h279 : ret <= 8'h33;
  11'h27a : ret <= 8'ha;
  11'h27b : ret <= 8'h32;
  11'h27c : ret <= 8'ha;
  11'h27d : ret <= 8'h31;
  11'h27e : ret <= 8'hd;
  11'h27f : ret <= 8'h22;
  11'h280 : ret <= 8'hb;
  11'h281 : ret <= 8'h23;
  11'h282 : ret <= 8'hb;
  11'h283 : ret <= 8'h24;
  11'h284 : ret <= 8'hb;
  11'h285 : ret <= 8'h25;
  11'h286 : ret <= 8'hb;
  11'h287 : ret <= 8'h26;
  11'h288 : ret <= 8'hb;
  11'h289 : ret <= 8'h27;
  11'h28a : ret <= 8'hb;
  11'h28b : ret <= 8'h28;
  11'h28c : ret <= 8'hb;
  11'h28d : ret <= 8'h21;
  11'h28e : ret <= 8'hb;
  11'h28f : ret <= 8'h14;
  11'h290 : ret <= 8'h3c;
  11'h291 : ret <= 8'h10;
  11'h292 : ret <= 8'h3b;
  11'h293 : ret <= 8'h10;
  11'h294 : ret <= 8'h7b;
  11'h295 : ret <= 8'hac;
  11'h296 : ret <= 8'h3b;
  11'h297 : ret <= 8'h11;
  11'h298 : ret <= 8'h7b;
  11'h299 : ret <= 8'hac;
  11'h29a : ret <= 8'h3b;
  11'h29b : ret <= 8'h1e;
  11'h29c : ret <= 8'h7b;
  11'h29d : ret <= 8'hac;
  11'h29e : ret <= 8'h3b;
  11'h29f : ret <= 8'h1c;
  11'h2a0 : ret <= 8'h7b;
  11'h2a1 : ret <= 8'hc;
  11'h2a2 : ret <= 8'h21;
  11'h2a3 : ret <= 8'h32;
  11'h2a4 : ret <= 8'ha;
  11'h2a5 : ret <= 8'h31;
  11'h2a6 : ret <= 8'h10;
  11'h2a7 : ret <= 8'h33;
  11'h2a8 : ret <= 8'h11;
  11'h2a9 : ret <= 8'h3c;
  11'h2aa : ret <= 8'h22;
  11'h2ab : ret <= 8'hbc;
  11'h2ac : ret <= 8'h34;
  11'h2ad : ret <= 8'h14;
  11'h2ae : ret <= 8'h3c;
  11'h2af : ret <= 8'h10;
  11'h2b0 : ret <= 8'h3b;
  11'h2b1 : ret <= 8'h10;
  11'h2b2 : ret <= 8'h7b;
  11'h2b3 : ret <= 8'hac;
  11'h2b4 : ret <= 8'h3b;
  11'h2b5 : ret <= 8'h12;
  11'h2b6 : ret <= 8'h7b;
  11'h2b7 : ret <= 8'hac;
  11'h2b8 : ret <= 8'h3b;
  11'h2b9 : ret <= 8'h1d;
  11'h2ba : ret <= 8'h7b;
  11'h2bb : ret <= 8'hac;
  11'h2bc : ret <= 8'h3b;
  11'h2bd : ret <= 8'h19;
  11'h2be : ret <= 8'h7b;
  11'h2bf : ret <= 8'h35;
  11'h2c0 : ret <= 8'h14;
  11'h2c1 : ret <= 8'h3c;
  11'h2c2 : ret <= 8'h10;
  11'h2c3 : ret <= 8'h3b;
  11'h2c4 : ret <= 8'h10;
  11'h2c5 : ret <= 8'h7b;
  11'h2c6 : ret <= 8'hac;
  11'h2c7 : ret <= 8'h3b;
  11'h2c8 : ret <= 8'h12;
  11'h2c9 : ret <= 8'h7b;
  11'h2ca : ret <= 8'hac;
  11'h2cb : ret <= 8'h3b;
  11'h2cc : ret <= 8'h1f;
  11'h2cd : ret <= 8'h7b;
  11'h2ce : ret <= 8'hac;
  11'h2cf : ret <= 8'h3b;
  11'h2d0 : ret <= 8'h14;
  11'h2d1 : ret <= 8'h7b;
  11'h2d2 : ret <= 8'h36;
  11'h2d3 : ret <= 8'hb;
  11'h2d4 : ret <= 8'h2d;
  11'h2d5 : ret <= 8'h37;
  11'h2d6 : ret <= 8'ha;
  11'h2d7 : ret <= 8'h16;
  11'h2d8 : ret <= 8'h3d;
  11'h2d9 : ret <= 8'h23;
  11'h2da : ret <= 8'hc4;
  11'h2db : ret <= 8'h26;
  11'h2dc : ret <= 8'h9;
  11'h2dd : ret <= 8'h21;
  11'h2de : ret <= 8'h43;
  11'h2df : ret <= 8'h3b;
  11'h2e0 : ret <= 8'hf0;
  11'h2e1 : ret <= 8'hb;
  11'h2e2 : ret <= 8'h11;
  11'h2e3 : ret <= 8'h3c;
  11'h2e4 : ret <= 8'h21;
  11'h2e5 : ret <= 8'h42;
  11'h2e6 : ret <= 8'h53;
  11'h2e7 : ret <= 8'h5c;
  11'h2e8 : ret <= 8'h3c;
  11'h2e9 : ret <= 8'hfc;
  11'h2ea : ret <= 8'h38;
  11'h2eb : ret <= 8'ha;
  11'h2ec : ret <= 8'hec;
  11'h2ed : ret <= 8'h28;
  11'h2ee : ret <= 8'heb;
  11'h2ef : ret <= 8'h11;
  11'h2f0 : ret <= 8'h43;
  11'h2f1 : ret <= 8'h33;
  11'h2f2 : ret <= 8'h25;
  11'h2f3 : ret <= 8'h8;
  11'h2f4 : ret <= 8'h27;
  11'h2f5 : ret <= 8'h3d;
  11'h2f6 : ret <= 8'ha;
  11'h2f7 : ret <= 8'h38;
  11'h2f8 : ret <= 8'ha;
  11'h2f9 : ret <= 8'h37;
  11'h2fa : ret <= 8'ha;
  11'h2fb : ret <= 8'h36;
  11'h2fc : ret <= 8'ha;
  11'h2fd : ret <= 8'h35;
  11'h2fe : ret <= 8'ha;
  11'h2ff : ret <= 8'h34;
  11'h300 : ret <= 8'ha;
  11'h301 : ret <= 8'h33;
  11'h302 : ret <= 8'ha;
  11'h303 : ret <= 8'h32;
  11'h304 : ret <= 8'hd;
  11'h305 : ret <= 8'h21;
  11'h306 : ret <= 8'hb;
  11'h307 : ret <= 8'h22;
  11'h308 : ret <= 8'hb;
  11'h309 : ret <= 8'h23;
  11'h30a : ret <= 8'hb;
  11'h30b : ret <= 8'h24;
  11'h30c : ret <= 8'hb;
  11'h30d : ret <= 8'h25;
  11'h30e : ret <= 8'hb;
  11'h30f : ret <= 8'h26;
  11'h310 : ret <= 8'hb;
  11'h311 : ret <= 8'h14;
  11'h312 : ret <= 8'h3c;
  11'h313 : ret <= 8'h10;
  11'h314 : ret <= 8'h3b;
  11'h315 : ret <= 8'h10;
  11'h316 : ret <= 8'h7b;
  11'h317 : ret <= 8'hac;
  11'h318 : ret <= 8'h3b;
  11'h319 : ret <= 8'h13;
  11'h31a : ret <= 8'h7b;
  11'h31b : ret <= 8'hac;
  11'h31c : ret <= 8'h3b;
  11'h31d : ret <= 8'h14;
  11'h31e : ret <= 8'h7b;
  11'h31f : ret <= 8'hac;
  11'h320 : ret <= 8'h3b;
  11'h321 : ret <= 8'h1c;
  11'h322 : ret <= 8'h7b;
  11'h323 : ret <= 8'h33;
  11'h324 : ret <= 8'h14;
  11'h325 : ret <= 8'h3c;
  11'h326 : ret <= 8'h10;
  11'h327 : ret <= 8'h3b;
  11'h328 : ret <= 8'h10;
  11'h329 : ret <= 8'h7b;
  11'h32a : ret <= 8'hac;
  11'h32b : ret <= 8'h3b;
  11'h32c : ret <= 8'h13;
  11'h32d : ret <= 8'h7b;
  11'h32e : ret <= 8'hac;
  11'h32f : ret <= 8'h3b;
  11'h330 : ret <= 8'h16;
  11'h331 : ret <= 8'h7b;
  11'h332 : ret <= 8'hac;
  11'h333 : ret <= 8'h3b;
  11'h334 : ret <= 8'h14;
  11'h335 : ret <= 8'h7b;
  11'h336 : ret <= 8'h34;
  11'h337 : ret <= 8'h11;
  11'h338 : ret <= 8'h35;
  11'h339 : ret <= 8'h14;
  11'h33a : ret <= 8'h3c;
  11'h33b : ret <= 8'h10;
  11'h33c : ret <= 8'h3b;
  11'h33d : ret <= 8'h10;
  11'h33e : ret <= 8'h7b;
  11'h33f : ret <= 8'hac;
  11'h340 : ret <= 8'h3b;
  11'h341 : ret <= 8'h10;
  11'h342 : ret <= 8'h7b;
  11'h343 : ret <= 8'hac;
  11'h344 : ret <= 8'h3b;
  11'h345 : ret <= 8'h18;
  11'h346 : ret <= 8'h7b;
  11'h347 : ret <= 8'hac;
  11'h348 : ret <= 8'h3b;
  11'h349 : ret <= 8'h17;
  11'h34a : ret <= 8'h7b;
  11'h34b : ret <= 8'h36;
  11'h34c : ret <= 8'h10;
  11'h34d : ret <= 8'hc2;
  11'h34e : ret <= 8'h24;
  11'h34f : ret <= 8'h9;
  11'h350 : ret <= 8'hf1;
  11'h351 : ret <= 8'h3c;
  11'h352 : ret <= 8'h21;
  11'h353 : ret <= 8'hb;
  11'h354 : ret <= 8'hb;
  11'h355 : ret <= 8'h2c;
  11'h356 : ret <= 8'h31;
  11'h357 : ret <= 8'ha;
  11'h358 : ret <= 8'h26;
  11'h359 : ret <= 8'hc;
  11'h35a : ret <= 8'ha;
  11'h35b : ret <= 8'h31;
  11'h35c : ret <= 8'h21;
  11'h35d : ret <= 8'h45;
  11'h35e : ret <= 8'h31;
  11'h35f : ret <= 8'h22;
  11'h360 : ret <= 8'h55;
  11'h361 : ret <= 8'h32;
  11'h362 : ret <= 8'h23;
  11'h363 : ret <= 8'h8;
  11'h364 : ret <= 8'ha;
  11'h365 : ret <= 8'h36;
  11'h366 : ret <= 8'ha;
  11'h367 : ret <= 8'h35;
  11'h368 : ret <= 8'ha;
  11'h369 : ret <= 8'h34;
  11'h36a : ret <= 8'ha;
  11'h36b : ret <= 8'h33;
  11'h36c : ret <= 8'ha;
  11'h36d : ret <= 8'h32;
  11'h36e : ret <= 8'ha;
  11'h36f : ret <= 8'h31;
  11'h370 : ret <= 8'hd;
  11'h371 : ret <= 8'h22;
  11'h372 : ret <= 8'hb;
  11'h373 : ret <= 8'h21;
  11'h374 : ret <= 8'hb;
  11'h375 : ret <= 8'h14;
  11'h376 : ret <= 8'h3c;
  11'h377 : ret <= 8'h10;
  11'h378 : ret <= 8'h3b;
  11'h379 : ret <= 8'h10;
  11'h37a : ret <= 8'h7b;
  11'h37b : ret <= 8'hac;
  11'h37c : ret <= 8'h3b;
  11'h37d : ret <= 8'h11;
  11'h37e : ret <= 8'h7b;
  11'h37f : ret <= 8'hac;
  11'h380 : ret <= 8'h3b;
  11'h381 : ret <= 8'h1e;
  11'h382 : ret <= 8'h7b;
  11'h383 : ret <= 8'hac;
  11'h384 : ret <= 8'h3b;
  11'h385 : ret <= 8'h1c;
  11'h386 : ret <= 8'h7b;
  11'h387 : ret <= 8'hc;
  11'h388 : ret <= 8'hb;
  11'h389 : ret <= 8'h21;
  11'h38a : ret <= 8'h32;
  11'h38b : ret <= 8'ha;
  11'h38c : ret <= 8'ha;
  11'h38d : ret <= 8'h31;
  11'h38e : ret <= 8'h14;
  11'h38f : ret <= 8'h3c;
  11'h390 : ret <= 8'h10;
  11'h391 : ret <= 8'h3b;
  11'h392 : ret <= 8'h10;
  11'h393 : ret <= 8'h7b;
  11'h394 : ret <= 8'hac;
  11'h395 : ret <= 8'h3b;
  11'h396 : ret <= 8'h13;
  11'h397 : ret <= 8'h7b;
  11'h398 : ret <= 8'hac;
  11'h399 : ret <= 8'h3b;
  11'h39a : ret <= 8'h10;
  11'h39b : ret <= 8'h7b;
  11'h39c : ret <= 8'hac;
  11'h39d : ret <= 8'h3b;
  11'h39e : ret <= 8'h15;
  11'h39f : ret <= 8'h7b;
  11'h3a0 : ret <= 8'hc;
  11'h3a1 : ret <= 8'ha;
  11'h3a2 : ret <= 8'h32;
  11'h3a3 : ret <= 8'hd;
  11'h3a4 : ret <= 8'h10;
  11'h3a5 : ret <= 8'hc1;
  11'h3a6 : ret <= 8'h14;
  11'h3a7 : ret <= 8'h3c;
  11'h3a8 : ret <= 8'h10;
  11'h3a9 : ret <= 8'h3b;
  11'h3aa : ret <= 8'h10;
  11'h3ab : ret <= 8'h7b;
  11'h3ac : ret <= 8'hac;
  11'h3ad : ret <= 8'h3b;
  11'h3ae : ret <= 8'h14;
  11'h3af : ret <= 8'h7b;
  11'h3b0 : ret <= 8'hac;
  11'h3b1 : ret <= 8'h3b;
  11'h3b2 : ret <= 8'h15;
  11'h3b3 : ret <= 8'h7b;
  11'h3b4 : ret <= 8'hac;
  11'h3b5 : ret <= 8'h3b;
  11'h3b6 : ret <= 8'h14;
  11'h3b7 : ret <= 8'h7b;
  11'h3b8 : ret <= 8'h9;
  11'h3b9 : ret <= 8'h21;
  11'h3ba : ret <= 8'hb;
  11'h3bb : ret <= 8'h22;
  11'h3bc : ret <= 8'hb;
  11'h3bd : ret <= 8'h23;
  11'h3be : ret <= 8'hb;
  11'h3bf : ret <= 8'h24;
  11'h3c0 : ret <= 8'hb;
  11'h3c1 : ret <= 8'h25;
  11'h3c2 : ret <= 8'hb;
  11'h3c3 : ret <= 8'h26;
  11'h3c4 : ret <= 8'hb;
  11'h3c5 : ret <= 8'h27;
  11'h3c6 : ret <= 8'hb;
  11'h3c7 : ret <= 8'hb;
  11'h3c8 : ret <= 8'h22;
  11'h3c9 : ret <= 8'h33;
  11'h3ca : ret <= 8'ha;
  11'h3cb : ret <= 8'h14;
  11'h3cc : ret <= 8'h3c;
  11'h3cd : ret <= 8'h10;
  11'h3ce : ret <= 8'h3b;
  11'h3cf : ret <= 8'h10;
  11'h3d0 : ret <= 8'h7b;
  11'h3d1 : ret <= 8'hac;
  11'h3d2 : ret <= 8'h3b;
  11'h3d3 : ret <= 8'h14;
  11'h3d4 : ret <= 8'h7b;
  11'h3d5 : ret <= 8'hac;
  11'h3d6 : ret <= 8'h3b;
  11'h3d7 : ret <= 8'h11;
  11'h3d8 : ret <= 8'h7b;
  11'h3d9 : ret <= 8'hac;
  11'h3da : ret <= 8'h3b;
  11'h3db : ret <= 8'h1b;
  11'h3dc : ret <= 8'h7b;
  11'h3dd : ret <= 8'h36;
  11'h3de : ret <= 8'hb;
  11'h3df : ret <= 8'h14;
  11'h3e0 : ret <= 8'h3c;
  11'h3e1 : ret <= 8'h10;
  11'h3e2 : ret <= 8'h3b;
  11'h3e3 : ret <= 8'h10;
  11'h3e4 : ret <= 8'h7b;
  11'h3e5 : ret <= 8'hac;
  11'h3e6 : ret <= 8'h3b;
  11'h3e7 : ret <= 8'h10;
  11'h3e8 : ret <= 8'h7b;
  11'h3e9 : ret <= 8'hac;
  11'h3ea : ret <= 8'h3b;
  11'h3eb : ret <= 8'h10;
  11'h3ec : ret <= 8'h7b;
  11'h3ed : ret <= 8'hac;
  11'h3ee : ret <= 8'h3b;
  11'h3ef : ret <= 8'h1a;
  11'h3f0 : ret <= 8'h7b;
  11'h3f1 : ret <= 8'h34;
  11'h3f2 : ret <= 8'ha;
  11'h3f3 : ret <= 8'hb;
  11'h3f4 : ret <= 8'h14;
  11'h3f5 : ret <= 8'h3c;
  11'h3f6 : ret <= 8'h10;
  11'h3f7 : ret <= 8'h3b;
  11'h3f8 : ret <= 8'h10;
  11'h3f9 : ret <= 8'h7b;
  11'h3fa : ret <= 8'hac;
  11'h3fb : ret <= 8'h3b;
  11'h3fc : ret <= 8'h10;
  11'h3fd : ret <= 8'h7b;
  11'h3fe : ret <= 8'hac;
  11'h3ff : ret <= 8'h3b;
  11'h400 : ret <= 8'h13;
  11'h401 : ret <= 8'h7b;
  11'h402 : ret <= 8'hac;
  11'h403 : ret <= 8'h3b;
  11'h404 : ret <= 8'h10;
  11'h405 : ret <= 8'h7b;
  11'h406 : ret <= 8'h35;
  11'h407 : ret <= 8'ha;
  11'h408 : ret <= 8'h14;
  11'h409 : ret <= 8'h3c;
  11'h40a : ret <= 8'h10;
  11'h40b : ret <= 8'h3b;
  11'h40c : ret <= 8'h10;
  11'h40d : ret <= 8'h7b;
  11'h40e : ret <= 8'hac;
  11'h40f : ret <= 8'h3b;
  11'h410 : ret <= 8'h11;
  11'h411 : ret <= 8'h7b;
  11'h412 : ret <= 8'hac;
  11'h413 : ret <= 8'h3b;
  11'h414 : ret <= 8'h13;
  11'h415 : ret <= 8'h7b;
  11'h416 : ret <= 8'hac;
  11'h417 : ret <= 8'h3b;
  11'h418 : ret <= 8'h1c;
  11'h419 : ret <= 8'h7b;
  11'h41a : ret <= 8'h37;
  11'h41b : ret <= 8'hb;
  11'h41c : ret <= 8'h24;
  11'h41d : ret <= 8'h32;
  11'h41e : ret <= 8'ha;
  11'h41f : ret <= 8'h27;
  11'h420 : ret <= 8'hc;
  11'h421 : ret <= 8'h22;
  11'h422 : ret <= 8'h45;
  11'h423 : ret <= 8'he3;
  11'h424 : ret <= 8'h11;
  11'h425 : ret <= 8'h43;
  11'h426 : ret <= 8'h33;
  11'h427 : ret <= 8'h10;
  11'h428 : ret <= 8'hc1;
  11'h429 : ret <= 8'h26;
  11'h42a : ret <= 8'h1;
  11'h42b : ret <= 8'h9;
  11'h42c : ret <= 8'h10;
  11'h42d : ret <= 8'he3;
  11'h42e : ret <= 8'ha;
  11'h42f : ret <= 8'h37;
  11'h430 : ret <= 8'ha;
  11'h431 : ret <= 8'h36;
  11'h432 : ret <= 8'ha;
  11'h433 : ret <= 8'h35;
  11'h434 : ret <= 8'ha;
  11'h435 : ret <= 8'h34;
  11'h436 : ret <= 8'ha;
  11'h437 : ret <= 8'h33;
  11'h438 : ret <= 8'ha;
  11'h439 : ret <= 8'h32;
  11'h43a : ret <= 8'hb;
  11'h43b : ret <= 8'h22;
  11'h43c : ret <= 8'h31;
  11'h43d : ret <= 8'ha;
  11'h43e : ret <= 8'h14;
  11'h43f : ret <= 8'h3c;
  11'h440 : ret <= 8'h10;
  11'h441 : ret <= 8'h3b;
  11'h442 : ret <= 8'h10;
  11'h443 : ret <= 8'h7b;
  11'h444 : ret <= 8'hac;
  11'h445 : ret <= 8'h3b;
  11'h446 : ret <= 8'h12;
  11'h447 : ret <= 8'h7b;
  11'h448 : ret <= 8'hac;
  11'h449 : ret <= 8'h3b;
  11'h44a : ret <= 8'h17;
  11'h44b : ret <= 8'h7b;
  11'h44c : ret <= 8'hac;
  11'h44d : ret <= 8'h3b;
  11'h44e : ret <= 8'h1f;
  11'h44f : ret <= 8'h7b;
  11'h450 : ret <= 8'hc;
  11'h451 : ret <= 8'ha;
  11'h452 : ret <= 8'h31;
  11'h453 : ret <= 8'hd;
  11'h454 : ret <= 8'h14;
  11'h455 : ret <= 8'h3c;
  11'h456 : ret <= 8'h10;
  11'h457 : ret <= 8'h3b;
  11'h458 : ret <= 8'h10;
  11'h459 : ret <= 8'h7b;
  11'h45a : ret <= 8'hac;
  11'h45b : ret <= 8'h3b;
  11'h45c : ret <= 8'h10;
  11'h45d : ret <= 8'h7b;
  11'h45e : ret <= 8'hac;
  11'h45f : ret <= 8'h3b;
  11'h460 : ret <= 8'h13;
  11'h461 : ret <= 8'h7b;
  11'h462 : ret <= 8'hac;
  11'h463 : ret <= 8'h3b;
  11'h464 : ret <= 8'h10;
  11'h465 : ret <= 8'h7b;
  11'h466 : ret <= 8'he2;
  11'h467 : ret <= 8'h11;
  11'h468 : ret <= 8'h42;
  11'h469 : ret <= 8'hec;
  11'h46a : ret <= 8'h10;
  11'h46b : ret <= 8'hec;
  11'h46c : ret <= 8'hd;
  11'h46d : ret <= 8'h22;
  11'h46e : ret <= 8'hb;
  11'h46f : ret <= 8'h14;
  11'h470 : ret <= 8'h3c;
  11'h471 : ret <= 8'h10;
  11'h472 : ret <= 8'h3b;
  11'h473 : ret <= 8'h10;
  11'h474 : ret <= 8'h7b;
  11'h475 : ret <= 8'hac;
  11'h476 : ret <= 8'h3b;
  11'h477 : ret <= 8'h10;
  11'h478 : ret <= 8'h7b;
  11'h479 : ret <= 8'hac;
  11'h47a : ret <= 8'h3b;
  11'h47b : ret <= 8'h16;
  11'h47c : ret <= 8'h7b;
  11'h47d : ret <= 8'hac;
  11'h47e : ret <= 8'h3b;
  11'h47f : ret <= 8'h14;
  11'h480 : ret <= 8'h7b;
  11'h481 : ret <= 8'h4f;
  11'h482 : ret <= 8'h32;
  11'h483 : ret <= 8'h14;
  11'h484 : ret <= 8'h3c;
  11'h485 : ret <= 8'h10;
  11'h486 : ret <= 8'h3b;
  11'h487 : ret <= 8'h10;
  11'h488 : ret <= 8'h7b;
  11'h489 : ret <= 8'hac;
  11'h48a : ret <= 8'h3b;
  11'h48b : ret <= 8'h13;
  11'h48c : ret <= 8'h7b;
  11'h48d : ret <= 8'hac;
  11'h48e : ret <= 8'h3b;
  11'h48f : ret <= 8'h1a;
  11'h490 : ret <= 8'h7b;
  11'h491 : ret <= 8'hac;
  11'h492 : ret <= 8'h3b;
  11'h493 : ret <= 8'h14;
  11'h494 : ret <= 8'h7b;
  11'h495 : ret <= 8'hc;
  11'h496 : ret <= 8'h21;
  11'h497 : ret <= 8'hb;
  11'h498 : ret <= 8'hb;
  11'h499 : ret <= 8'h22;
  11'h49a : ret <= 8'h31;
  11'h49b : ret <= 8'ha;
  11'h49c : ret <= 8'h14;
  11'h49d : ret <= 8'h3c;
  11'h49e : ret <= 8'h10;
  11'h49f : ret <= 8'h3b;
  11'h4a0 : ret <= 8'h10;
  11'h4a1 : ret <= 8'h7b;
  11'h4a2 : ret <= 8'hac;
  11'h4a3 : ret <= 8'h3b;
  11'h4a4 : ret <= 8'h13;
  11'h4a5 : ret <= 8'h7b;
  11'h4a6 : ret <= 8'hac;
  11'h4a7 : ret <= 8'h3b;
  11'h4a8 : ret <= 8'h17;
  11'h4a9 : ret <= 8'h7b;
  11'h4aa : ret <= 8'hac;
  11'h4ab : ret <= 8'h3b;
  11'h4ac : ret <= 8'h11;
  11'h4ad : ret <= 8'h7b;
  11'h4ae : ret <= 8'hc;
  11'h4af : ret <= 8'ha;
  11'h4b0 : ret <= 8'h31;
  11'h4b1 : ret <= 8'ha;
  11'h4b2 : ret <= 8'h32;
  11'h4b3 : ret <= 8'hd;
  11'h4b4 : ret <= 8'h0;
  default: ret <= 8'h0;
endcase
endmodule

module rom2_wide(input clk, input enable ,input [10:0] addr, output [15:0] data_out);
rom2 rom2_low(clk, enable, addr, data_out[7:0]);
rom2 rom2_high(clk, enable, addr+11'h1, data_out[15:8]);
endmodule

