module reflet_bootloader16_rom(input clk, input enable, input [14-1:0] addr, output [16-1:0] data);
    reg [16-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            14'h3E80 : data_reg <= 16'h1220;
            14'h3E81 : data_reg <= 16'h1124;
            14'h3E82 : data_reg <= 16'h1B0D;
            14'h3E83 : data_reg <= 16'h1C28;
            14'h3E84 : data_reg <= 16'h8C22;
            14'h3E85 : data_reg <= 16'h9C6D;
            14'h3E86 : data_reg <= 16'h6D8C;
            14'h3E87 : data_reg <= 16'h221D;
            14'h3E88 : data_reg <= 16'h001C;
            14'h3E89 : data_reg <= 16'h3C22;
            14'h3E8A : data_reg <= 16'h1E3E;
            14'h3E8B : data_reg <= 16'h7F60;
            14'h3E8C : data_reg <= 16'h3C23;
            14'h3E8D : data_reg <= 16'h3EE5;
            14'h3E8E : data_reg <= 16'h1CD0;
            14'h3E8F : data_reg <= 16'h1D0B;
            14'h3E90 : data_reg <= 16'hD00C;
            14'h3E91 : data_reg <= 16'h2813;
            14'h3E92 : data_reg <= 16'h211C;
            14'h3E93 : data_reg <= 16'h6D8C;
            14'h3E94 : data_reg <= 16'h8C9C;
            14'h3E95 : data_reg <= 16'h1D6D;
            14'h3E96 : data_reg <= 16'h14D3;
            14'h3E97 : data_reg <= 16'h3321;
            14'h3E98 : data_reg <= 16'hD313;
            14'h3E99 : data_reg <= 16'h2F15;
            14'h3E9A : data_reg <= 16'h1333;
            14'h3E9B : data_reg <= 16'h1B0D;
            14'h3E9C : data_reg <= 16'h1C28;
            14'h3E9D : data_reg <= 16'h8C22;
            14'h3E9E : data_reg <= 16'h9C6D;
            14'h3E9F : data_reg <= 16'h6D8C;
            14'h3EA0 : data_reg <= 16'h221D;
            14'h3EA1 : data_reg <= 16'h001C;
            14'h3EA2 : data_reg <= 16'h3C22;
            14'h3EA3 : data_reg <= 16'h1E3E;
            14'h3EA4 : data_reg <= 16'h0063;
            14'h3EA5 : data_reg <= 16'h3C23;
            14'h3EA6 : data_reg <= 16'h3EE5;
            14'h3EA7 : data_reg <= 16'h1CD0;
            14'h3EA8 : data_reg <= 16'h1D0B;
            14'h3EA9 : data_reg <= 16'hC30C;
            14'h3EAA : data_reg <= 16'h2116;
            14'h3EAB : data_reg <= 16'h1333;
            14'h3EAC : data_reg <= 16'hC306;
            14'h3EAD : data_reg <= 16'h3321;
            14'h3EAE : data_reg <= 16'h2113;
            14'h3EAF : data_reg <= 16'h20C3;
            14'h3EB0 : data_reg <= 16'hE6A5;
            14'h3EB1 : data_reg <= 16'h1B0D;
            14'h3EB2 : data_reg <= 16'h1C28;
            14'h3EB3 : data_reg <= 16'h8C22;
            14'h3EB4 : data_reg <= 16'h9C6D;
            14'h3EB5 : data_reg <= 16'h6D8C;
            14'h3EB6 : data_reg <= 16'h221D;
            14'h3EB7 : data_reg <= 16'h001C;
            14'h3EB8 : data_reg <= 16'h3C22;
            14'h3EB9 : data_reg <= 16'h1E3E;
            14'h3EBA : data_reg <= 16'h7DA8;
            14'h3EBB : data_reg <= 16'h3C23;
            14'h3EBC : data_reg <= 16'h3EE5;
            14'h3EBD : data_reg <= 16'h1CD0;
            14'h3EBE : data_reg <= 16'h1D0B;
            14'h3EBF : data_reg <= 16'hE00C;
            14'h3EC0 : data_reg <= 16'h3321;
            14'h3EC1 : data_reg <= 16'h2113;
            14'h3EC2 : data_reg <= 16'h22C3;
            14'h3EC3 : data_reg <= 16'h1333;
            14'h3EC4 : data_reg <= 16'hC304;
            14'h3EC5 : data_reg <= 16'h1B0D;
            14'h3EC6 : data_reg <= 16'h1C28;
            14'h3EC7 : data_reg <= 16'h8C22;
            14'h3EC8 : data_reg <= 16'h9C6D;
            14'h3EC9 : data_reg <= 16'h6D8C;
            14'h3ECA : data_reg <= 16'h221D;
            14'h3ECB : data_reg <= 16'h001C;
            14'h3ECC : data_reg <= 16'h3C22;
            14'h3ECD : data_reg <= 16'h1E3E;
            14'h3ECE : data_reg <= 16'h7DD3;
            14'h3ECF : data_reg <= 16'h3C23;
            14'h3ED0 : data_reg <= 16'h3EE5;
            14'h3ED1 : data_reg <= 16'h1CD0;
            14'h3ED2 : data_reg <= 16'h1D0B;
            14'h3ED3 : data_reg <= 16'h1E0C;
            14'h3ED4 : data_reg <= 16'h3321;
            14'h3ED5 : data_reg <= 16'h2113;
            14'h3ED6 : data_reg <= 16'h21C3;
            14'h3ED7 : data_reg <= 16'h1333;
            14'h3ED8 : data_reg <= 16'h1B0D;
            14'h3ED9 : data_reg <= 16'h1C28;
            14'h3EDA : data_reg <= 16'h8C22;
            14'h3EDB : data_reg <= 16'h9C6D;
            14'h3EDC : data_reg <= 16'h6D8C;
            14'h3EDD : data_reg <= 16'h221D;
            14'h3EDE : data_reg <= 16'h001C;
            14'h3EDF : data_reg <= 16'h3C22;
            14'h3EE0 : data_reg <= 16'h1E3E;
            14'h3EE1 : data_reg <= 16'h00FF;
            14'h3EE2 : data_reg <= 16'h3C23;
            14'h3EE3 : data_reg <= 16'h3EE5;
            14'h3EE4 : data_reg <= 16'h1CD0;
            14'h3EE5 : data_reg <= 16'h1D0B;
            14'h3EE6 : data_reg <= 16'hC30C;
            14'h3EE7 : data_reg <= 16'h3321;
            14'h3EE8 : data_reg <= 16'h0513;
            14'h3EE9 : data_reg <= 16'h0DC3;
            14'h3EEA : data_reg <= 16'h281B;
            14'h3EEB : data_reg <= 16'h221C;
            14'h3EEC : data_reg <= 16'h6D8C;
            14'h3EED : data_reg <= 16'h8C9C;
            14'h3EEE : data_reg <= 16'h1D6D;
            14'h3EEF : data_reg <= 16'h1C22;
            14'h3EF0 : data_reg <= 16'h3C22;
            14'h3EF1 : data_reg <= 16'h1E3E;
            14'h3EF2 : data_reg <= 16'h7F62;
            14'h3EF3 : data_reg <= 16'h3C23;
            14'h3EF4 : data_reg <= 16'h3EE5;
            14'h3EF5 : data_reg <= 16'h1CD0;
            14'h3EF6 : data_reg <= 16'h1D0B;
            14'h3EF7 : data_reg <= 16'h130C;
            14'h3EF8 : data_reg <= 16'h1B0D;
            14'h3EF9 : data_reg <= 16'h1C28;
            14'h3EFA : data_reg <= 16'h8C22;
            14'h3EFB : data_reg <= 16'h9C6D;
            14'h3EFC : data_reg <= 16'h6D8C;
            14'h3EFD : data_reg <= 16'hD31D;
            14'h3EFE : data_reg <= 16'h0B1C;
            14'h3EFF : data_reg <= 16'h0C1D;
            14'h3F00 : data_reg <= 16'h2A13;
            14'h3F01 : data_reg <= 16'h21C3;
            14'h3F02 : data_reg <= 16'h1333;
            14'h3F03 : data_reg <= 16'h1B0D;
            14'h3F04 : data_reg <= 16'h1C28;
            14'h3F05 : data_reg <= 16'h8C22;
            14'h3F06 : data_reg <= 16'h9C6D;
            14'h3F07 : data_reg <= 16'h6D8C;
            14'h3F08 : data_reg <= 16'h221D;
            14'h3F09 : data_reg <= 16'h001C;
            14'h3F0A : data_reg <= 16'h3C22;
            14'h3F0B : data_reg <= 16'h1E3E;
            14'h3F0C : data_reg <= 16'h0040;
            14'h3F0D : data_reg <= 16'h3C23;
            14'h3F0E : data_reg <= 16'h3EE5;
            14'h3F0F : data_reg <= 16'h1CD0;
            14'h3F10 : data_reg <= 16'h1D0B;
            14'h3F11 : data_reg <= 16'hC30C;
            14'h3F12 : data_reg <= 16'h3322;
            14'h3F13 : data_reg <= 16'h0D13;
            14'h3F14 : data_reg <= 16'h281B;
            14'h3F15 : data_reg <= 16'h221C;
            14'h3F16 : data_reg <= 16'h6D8C;
            14'h3F17 : data_reg <= 16'h8C9C;
            14'h3F18 : data_reg <= 16'h1D6D;
            14'h3F19 : data_reg <= 16'h1C22;
            14'h3F1A : data_reg <= 16'h3C22;
            14'h3F1B : data_reg <= 16'h1E3E;
            14'h3F1C : data_reg <= 16'h0190;
            14'h3F1D : data_reg <= 16'h3C23;
            14'h3F1E : data_reg <= 16'h3EE5;
            14'h3F1F : data_reg <= 16'h1CD0;
            14'h3F20 : data_reg <= 16'h1D0B;
            14'h3F21 : data_reg <= 16'h160C;
            14'h3F22 : data_reg <= 16'h0D11;
            14'h3F23 : data_reg <= 16'h281B;
            14'h3F24 : data_reg <= 16'h221C;
            14'h3F25 : data_reg <= 16'h6D8C;
            14'h3F26 : data_reg <= 16'h8C9C;
            14'h3F27 : data_reg <= 16'h1D6D;
            14'h3F28 : data_reg <= 16'h1C22;
            14'h3F29 : data_reg <= 16'h3C22;
            14'h3F2A : data_reg <= 16'h1E3E;
            14'h3F2B : data_reg <= 16'hFF19;
            14'h3F2C : data_reg <= 16'h3C23;
            14'h3F2D : data_reg <= 16'h3EE5;
            14'h3F2E : data_reg <= 16'h1CD0;
            14'h3F2F : data_reg <= 16'h1D0B;
            14'h3F30 : data_reg <= 16'h170C;
            14'h3F31 : data_reg <= 16'h1B0D;
            14'h3F32 : data_reg <= 16'h1C28;
            14'h3F33 : data_reg <= 16'h8C22;
            14'h3F34 : data_reg <= 16'h9C6D;
            14'h3F35 : data_reg <= 16'h6D8C;
            14'h3F36 : data_reg <= 16'h221D;
            14'h3F37 : data_reg <= 16'h001C;
            14'h3F38 : data_reg <= 16'h3C22;
            14'h3F39 : data_reg <= 16'h1E3E;
            14'h3F3A : data_reg <= 16'h7EE3;
            14'h3F3B : data_reg <= 16'h3C23;
            14'h3F3C : data_reg <= 16'h3EE5;
            14'h3F3D : data_reg <= 16'h1CD0;
            14'h3F3E : data_reg <= 16'h1D0B;
            14'h3F3F : data_reg <= 16'h180C;
            14'h3F40 : data_reg <= 16'h1B0D;
            14'h3F41 : data_reg <= 16'h1C28;
            14'h3F42 : data_reg <= 16'h8C22;
            14'h3F43 : data_reg <= 16'h9C6D;
            14'h3F44 : data_reg <= 16'h6D8C;
            14'h3F45 : data_reg <= 16'h221D;
            14'h3F46 : data_reg <= 16'h001C;
            14'h3F47 : data_reg <= 16'h3C22;
            14'h3F48 : data_reg <= 16'h1E3E;
            14'h3F49 : data_reg <= 16'h7F44;
            14'h3F4A : data_reg <= 16'h3C23;
            14'h3F4B : data_reg <= 16'h3EE5;
            14'h3F4C : data_reg <= 16'h1CD0;
            14'h3F4D : data_reg <= 16'h1D0B;
            14'h3F4E : data_reg <= 16'hEC0C;
            14'h3F4F : data_reg <= 16'h1B0D;
            14'h3F50 : data_reg <= 16'h1C28;
            14'h3F51 : data_reg <= 16'h8C22;
            14'h3F52 : data_reg <= 16'h9C6D;
            14'h3F53 : data_reg <= 16'h6D8C;
            14'h3F54 : data_reg <= 16'h221D;
            14'h3F55 : data_reg <= 16'h001C;
            14'h3F56 : data_reg <= 16'h3C22;
            14'h3F57 : data_reg <= 16'h1E3E;
            14'h3F58 : data_reg <= 16'h7F50;
            14'h3F59 : data_reg <= 16'h3C23;
            14'h3F5A : data_reg <= 16'h3EE5;
            14'h3F5B : data_reg <= 16'h1CD0;
            14'h3F5C : data_reg <= 16'h1D0B;
            14'h3F5D : data_reg <= 16'hED0C;
            14'h3F5E : data_reg <= 16'h5D26;
            14'h3F5F : data_reg <= 16'h0D1D;
            14'h3F60 : data_reg <= 16'h281B;
            14'h3F61 : data_reg <= 16'h221C;
            14'h3F62 : data_reg <= 16'h6D8C;
            14'h3F63 : data_reg <= 16'h8C9C;
            14'h3F64 : data_reg <= 16'h1D6D;
            14'h3F65 : data_reg <= 16'h1C22;
            14'h3F66 : data_reg <= 16'h3C22;
            14'h3F67 : data_reg <= 16'h1E3E;
            14'h3F68 : data_reg <= 16'h7EDC;
            14'h3F69 : data_reg <= 16'h3C23;
            14'h3F6A : data_reg <= 16'h3EE5;
            14'h3F6B : data_reg <= 16'h1CD0;
            14'h3F6C : data_reg <= 16'h1D0B;
            14'h3F6D : data_reg <= 16'h1A0C;
            14'h3F6E : data_reg <= 16'h2000;
            14'h3F6F : data_reg <= 16'h08A1;
            14'h3F70 : data_reg <= 16'h0AE0;
            14'h3F71 : data_reg <= 16'h281E;
            14'h3F72 : data_reg <= 16'h211C;
            14'h3F73 : data_reg <= 16'h6D8C;
            14'h3F74 : data_reg <= 16'h8C9C;
            14'h3F75 : data_reg <= 16'h1D6D;
            14'h3F76 : data_reg <= 16'h1B0D;
            14'h3F77 : data_reg <= 16'h1C28;
            14'h3F78 : data_reg <= 16'h8C22;
            14'h3F79 : data_reg <= 16'h9C6D;
            14'h3F7A : data_reg <= 16'h6D8C;
            14'h3F7B : data_reg <= 16'h221D;
            14'h3F7C : data_reg <= 16'h001C;
            14'h3F7D : data_reg <= 16'h3C22;
            14'h3F7E : data_reg <= 16'h1E3E;
            14'h3F7F : data_reg <= 16'hFF04;
            14'h3F80 : data_reg <= 16'h3C23;
            14'h3F81 : data_reg <= 16'h3EE5;
            14'h3F82 : data_reg <= 16'h1CD0;
            14'h3F83 : data_reg <= 16'h1D0B;
            14'h3F84 : data_reg <= 16'h110C;
            14'h3F85 : data_reg <= 16'hC120;
            14'h3F86 : data_reg <= 16'h3121;
            14'h3F87 : data_reg <= 16'h2011;
            14'h3F88 : data_reg <= 16'h21C1;
            14'h3F89 : data_reg <= 16'h1131;
            14'h3F8A : data_reg <= 16'hC120;
            14'h3F8B : data_reg <= 16'h3129;
            14'h3F8C : data_reg <= 16'h2011;
            14'h3F8D : data_reg <= 16'h21C1;
            14'h3F8E : data_reg <= 16'h1131;
            14'h3F8F : data_reg <= 16'hC120;
            14'h3F90 : data_reg <= 16'h3121;
            14'h3F91 : data_reg <= 16'h2011;
            14'h3F92 : data_reg <= 16'h21C1;
            14'h3F93 : data_reg <= 16'h1131;
            14'h3F94 : data_reg <= 16'hC120;
            14'h3F95 : data_reg <= 16'h3121;
            14'h3F96 : data_reg <= 16'h2011;
            14'h3F97 : data_reg <= 16'h21C1;
            14'h3F98 : data_reg <= 16'h1131;
            14'h3F99 : data_reg <= 16'hC120;
            14'h3F9A : data_reg <= 16'h1211;
            14'h3F9B : data_reg <= 16'h1413;
            14'h3F9C : data_reg <= 16'h1615;
            14'h3F9D : data_reg <= 16'h1817;
            14'h3F9E : data_reg <= 16'h1A19;
            14'h3F9F : data_reg <= 16'h1C1B;
            14'h3FA0 : data_reg <= 16'h1F1D;
            14'h3FA1 : data_reg <= 16'h1E24;
            14'h3FA2 : data_reg <= 16'h0614;
            14'h3FA3 : data_reg <= 16'h2011;
            14'h3FA4 : data_reg <= 16'hD7C3;
            14'h3FA5 : data_reg <= 16'h21C2;
            14'h3FA6 : data_reg <= 16'h1232;
            14'h3FA7 : data_reg <= 16'hEB04;
            14'h3FA8 : data_reg <= 16'h2015;
            14'h3FA9 : data_reg <= 16'h21C3;
            14'h3FAA : data_reg <= 16'h0119;
            14'h3FAB : data_reg <= 16'h39E5;
            14'h3FAC : data_reg <= 16'h11E5;
            14'h3FAD : data_reg <= 16'hEB05;
            14'h3FAE : data_reg <= 16'h7D00;
            14'h3FAF : data_reg <= 16'h8000;
            14'h3FB0 : data_reg <= 16'hFF00;
            14'h3FB1 : data_reg <= 16'hFF04;
            14'h3FB2 : data_reg <= 16'hFF08;
            14'h3FB3 : data_reg <= 16'hFF10;
            14'h3FB4 : data_reg <= 16'hFF13;
            14'h3FB5 : data_reg <= 16'hFF16;
            14'h3FB6 : data_reg <= 16'hFF1A;
            14'h3FB7 : data_reg <= 16'hFF1C;
            14'h3FB8 : data_reg <= 16'hFF1F;
            14'h3FB9 : data_reg <= 16'hFF21;
            14'h3FBA : data_reg <= 16'hFF22;
            default : data_reg <= 0;
        endcase
    assign data = ( enable ? data_reg : 0 );
endmodule
