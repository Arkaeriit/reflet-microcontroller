module rom07(input clk, input enable, input [8-1:0] addr, output [16-1:0] data);
    reg [16-1:0] data_reg;
    always @ (posedge clk)
        case(addr)
            8'h0 : data_reg <= 16'h5341;
            8'h1 : data_reg <= 16'h4D52;
            8'h2 : data_reg <= 16'h3C3C;
            8'h3 : data_reg <= 16'h3B2D;
            8'h4 : data_reg <= 16'h102C;
            8'h5 : data_reg <= 16'h123D;
            8'h6 : data_reg <= 16'h003C;
            8'h7 : data_reg <= 16'h0000;
            8'h8 : data_reg <= 16'h0000;
            8'h9 : data_reg <= 16'h4C12;
            8'hA : data_reg <= 16'h3E4E;
            8'hB : data_reg <= 16'h8000;
            8'hC : data_reg <= 16'h4C13;
            8'hD : data_reg <= 16'h4E08;
            8'hE : data_reg <= 16'h3CF0;
            8'hF : data_reg <= 16'h3D2B;
            8'h10 : data_reg <= 16'h3F2C;
            8'h11 : data_reg <= 16'h3C2C;
            8'h12 : data_reg <= 16'h3B2D;
            8'h13 : data_reg <= 16'h102C;
            8'h14 : data_reg <= 16'h123D;
            8'h15 : data_reg <= 16'h003C;
            8'h16 : data_reg <= 16'h0000;
            8'h17 : data_reg <= 16'h0000;
            8'h18 : data_reg <= 16'h4C12;
            8'h19 : data_reg <= 16'h3E4E;
            8'h1A : data_reg <= 16'h0173;
            8'h1B : data_reg <= 16'h4C13;
            8'h1C : data_reg <= 16'h4E08;
            8'h1D : data_reg <= 16'h3CF0;
            8'h1E : data_reg <= 16'h3D2B;
            8'h1F : data_reg <= 16'h3E2C;
            8'h20 : data_reg <= 16'h8000;
            8'h21 : data_reg <= 16'hFF00;
            8'h22 : data_reg <= 16'hFF04;
            8'h23 : data_reg <= 16'hFF08;
            8'h24 : data_reg <= 16'hFF10;
            8'h25 : data_reg <= 16'hFF13;
            8'h26 : data_reg <= 16'hFF16;
            8'h27 : data_reg <= 16'hFF1A;
            8'h28 : data_reg <= 16'hFF1C;
            8'h29 : data_reg <= 16'hFF1F;
            8'h2A : data_reg <= 16'hFF21;
            8'h2B : data_reg <= 16'hFF22;
            8'h2C : data_reg <= 16'h223C;
            8'h2D : data_reg <= 16'h2C0B;
            8'h2E : data_reg <= 16'h243C;
            8'h2F : data_reg <= 16'h2C0B;
            8'h30 : data_reg <= 16'h2D3C;
            8'h31 : data_reg <= 16'h2C3B;
            8'h32 : data_reg <= 16'h3D10;
            8'h33 : data_reg <= 16'h3C12;
            8'h34 : data_reg <= 16'h0000;
            8'h35 : data_reg <= 16'h0000;
            8'h36 : data_reg <= 16'h4C12;
            8'h37 : data_reg <= 16'h3E4E;
            8'h38 : data_reg <= 16'h004C;
            8'h39 : data_reg <= 16'h4C13;
            8'h3A : data_reg <= 16'h4E08;
            8'h3B : data_reg <= 16'h3CF0;
            8'h3C : data_reg <= 16'h3D2B;
            8'h3D : data_reg <= 16'hF02C;
            8'h3E : data_reg <= 16'h3203;
            8'h3F : data_reg <= 16'h2D3C;
            8'h40 : data_reg <= 16'h2C3B;
            8'h41 : data_reg <= 16'h3D10;
            8'h42 : data_reg <= 16'h3C12;
            8'h43 : data_reg <= 16'h0000;
            8'h44 : data_reg <= 16'h0000;
            8'h45 : data_reg <= 16'h4C12;
            8'h46 : data_reg <= 16'h3E4E;
            8'h47 : data_reg <= 16'h009A;
            8'h48 : data_reg <= 16'h4C13;
            8'h49 : data_reg <= 16'h4E08;
            8'h4A : data_reg <= 16'h3CF0;
            8'h4B : data_reg <= 16'h3D2B;
            8'h4C : data_reg <= 16'h342C;
            8'h4D : data_reg <= 16'h3CF2;
            8'h4E : data_reg <= 16'hCC10;
            8'h4F : data_reg <= 16'h0924;
            8'h50 : data_reg <= 16'h4211;
            8'h51 : data_reg <= 16'h213C;
            8'h52 : data_reg <= 16'h10EC;
            8'h53 : data_reg <= 16'h03E2;
            8'h54 : data_reg <= 16'h0A3C;
            8'h55 : data_reg <= 16'h2C34;
            8'h56 : data_reg <= 16'h0A3C;
            8'h57 : data_reg <= 16'h2C32;
            8'h58 : data_reg <= 16'h3C0D;
            8'h59 : data_reg <= 16'h0B21;
            8'h5A : data_reg <= 16'h1A2C;
            8'h5B : data_reg <= 16'h3C31;
            8'h5C : data_reg <= 16'h3B2D;
            8'h5D : data_reg <= 16'h102C;
            8'h5E : data_reg <= 16'h123D;
            8'h5F : data_reg <= 16'h003C;
            8'h60 : data_reg <= 16'h0000;
            8'h61 : data_reg <= 16'h0000;
            8'h62 : data_reg <= 16'h4C12;
            8'h63 : data_reg <= 16'h3E4E;
            8'h64 : data_reg <= 16'h0058;
            8'h65 : data_reg <= 16'h4C13;
            8'h66 : data_reg <= 16'h4E08;
            8'h67 : data_reg <= 16'h3CF0;
            8'h68 : data_reg <= 16'h3D2B;
            8'h69 : data_reg <= 16'h0C2C;
            8'h6A : data_reg <= 16'h311D;
            8'h6B : data_reg <= 16'h2D3C;
            8'h6C : data_reg <= 16'h2C3B;
            8'h6D : data_reg <= 16'h3D10;
            8'h6E : data_reg <= 16'h3C12;
            8'h6F : data_reg <= 16'h0000;
            8'h70 : data_reg <= 16'h0000;
            8'h71 : data_reg <= 16'h4C12;
            8'h72 : data_reg <= 16'h3E4E;
            8'h73 : data_reg <= 16'h0058;
            8'h74 : data_reg <= 16'h4C13;
            8'h75 : data_reg <= 16'h4E08;
            8'h76 : data_reg <= 16'h3CF0;
            8'h77 : data_reg <= 16'h3D2B;
            8'h78 : data_reg <= 16'h0C2C;
            8'h79 : data_reg <= 16'h0A3C;
            8'h7A : data_reg <= 16'h2C31;
            8'h7B : data_reg <= 16'h3C0D;
            8'h7C : data_reg <= 16'h0B22;
            8'h7D : data_reg <= 16'h3C2C;
            8'h7E : data_reg <= 16'h0B23;
            8'h7F : data_reg <= 16'h3C2C;
            8'h80 : data_reg <= 16'h3B2D;
            8'h81 : data_reg <= 16'h102C;
            8'h82 : data_reg <= 16'h123D;
            8'h83 : data_reg <= 16'h003C;
            8'h84 : data_reg <= 16'h0000;
            8'h85 : data_reg <= 16'h0000;
            8'h86 : data_reg <= 16'h4C12;
            8'h87 : data_reg <= 16'h3E4E;
            8'h88 : data_reg <= 16'h004C;
            8'h89 : data_reg <= 16'h4C13;
            8'h8A : data_reg <= 16'h4E08;
            8'h8B : data_reg <= 16'h3CF0;
            8'h8C : data_reg <= 16'h3D2B;
            8'h8D : data_reg <= 16'hF02C;
            8'h8E : data_reg <= 16'h1232;
            8'h8F : data_reg <= 16'h3242;
            8'h90 : data_reg <= 16'h2D3C;
            8'h91 : data_reg <= 16'h2C3B;
            8'h92 : data_reg <= 16'h3D10;
            8'h93 : data_reg <= 16'h3C12;
            8'h94 : data_reg <= 16'h0000;
            8'h95 : data_reg <= 16'h0000;
            8'h96 : data_reg <= 16'h4C12;
            8'h97 : data_reg <= 16'h3E4E;
            8'h98 : data_reg <= 16'h0141;
            8'h99 : data_reg <= 16'h4C13;
            8'h9A : data_reg <= 16'h4E08;
            8'h9B : data_reg <= 16'h3CF0;
            8'h9C : data_reg <= 16'h3D2B;
            8'h9D : data_reg <= 16'h332C;
            8'h9E : data_reg <= 16'h0311;
            8'h9F : data_reg <= 16'h03E2;
            8'hA0 : data_reg <= 16'h0331;
            8'hA1 : data_reg <= 16'h03F2;
            8'hA2 : data_reg <= 16'h23C1;
            8'hA3 : data_reg <= 16'h1109;
            8'hA4 : data_reg <= 16'h3242;
            8'hA5 : data_reg <= 16'hF203;
            8'hA6 : data_reg <= 16'h3103;
            8'hA7 : data_reg <= 16'h0A3C;
            8'hA8 : data_reg <= 16'h2C33;
            8'hA9 : data_reg <= 16'h0A3C;
            8'hAA : data_reg <= 16'h2C32;
            8'hAB : data_reg <= 16'h000D;
            8'hAC : data_reg <= 16'h0000;
            8'hAD : data_reg <= 16'h0000;
            8'hAE : data_reg <= 16'h0000;
            8'hAF : data_reg <= 16'h0000;
            8'hB0 : data_reg <= 16'h0000;
            8'hB1 : data_reg <= 16'h0000;
            8'hB2 : data_reg <= 16'h0000;
            8'hB3 : data_reg <= 16'h0000;
            8'hB4 : data_reg <= 16'h0000;
            8'hB5 : data_reg <= 16'h0000;
            8'hB6 : data_reg <= 16'h0000;
            8'hB7 : data_reg <= 16'h0000;
            8'hB8 : data_reg <= 16'h0000;
            8'hB9 : data_reg <= 16'h3C00;
            8'hBA : data_reg <= 16'h3B2D;
            8'hBB : data_reg <= 16'h102C;
            8'hBC : data_reg <= 16'h123D;
            8'hBD : data_reg <= 16'h003C;
            8'hBE : data_reg <= 16'h0000;
            8'hBF : data_reg <= 16'h0000;
            8'hC0 : data_reg <= 16'h4C12;
            8'hC1 : data_reg <= 16'h3E4E;
            8'hC2 : data_reg <= 16'h00F7;
            8'hC3 : data_reg <= 16'h4C13;
            8'hC4 : data_reg <= 16'h4E08;
            8'hC5 : data_reg <= 16'h3CF0;
            8'hC6 : data_reg <= 16'h3D2B;
            8'hC7 : data_reg <= 16'h0C2C;
            8'hC8 : data_reg <= 16'h2D3C;
            8'hC9 : data_reg <= 16'h2C3B;
            8'hCA : data_reg <= 16'h3D10;
            8'hCB : data_reg <= 16'h3C12;
            8'hCC : data_reg <= 16'h0000;
            8'hCD : data_reg <= 16'h0000;
            8'hCE : data_reg <= 16'h4C12;
            8'hCF : data_reg <= 16'h3E4E;
            8'hD0 : data_reg <= 16'h0058;
            8'hD1 : data_reg <= 16'h4C13;
            8'hD2 : data_reg <= 16'h4E08;
            8'hD3 : data_reg <= 16'h3CF0;
            8'hD4 : data_reg <= 16'h3D2B;
            8'hD5 : data_reg <= 16'h0C2C;
            8'hD6 : data_reg <= 16'h2D3C;
            8'hD7 : data_reg <= 16'h2C3B;
            8'hD8 : data_reg <= 16'h3D10;
            8'hD9 : data_reg <= 16'h3C12;
            8'hDA : data_reg <= 16'h0000;
            8'hDB : data_reg <= 16'h0000;
            8'hDC : data_reg <= 16'h4C12;
            8'hDD : data_reg <= 16'h3E4E;
            8'hDE : data_reg <= 16'h0173;
            8'hDF : data_reg <= 16'h4C13;
            8'hE0 : data_reg <= 16'h4E08;
            8'hE1 : data_reg <= 16'h3CF0;
            8'hE2 : data_reg <= 16'h3D2B;
            8'hE3 : data_reg <= 16'h3E2C;
            default : data_reg <= 0;
        endcase
    assign data = ( enable ? data_reg : 0 );
endmodule
